-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Oct 23 2024 20:10:58

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    start_stop : in std_logic;
    s2_phy : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    error_pin : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__53076\ : std_logic;
signal \N__53075\ : std_logic;
signal \N__53074\ : std_logic;
signal \N__53065\ : std_logic;
signal \N__53064\ : std_logic;
signal \N__53063\ : std_logic;
signal \N__53056\ : std_logic;
signal \N__53055\ : std_logic;
signal \N__53054\ : std_logic;
signal \N__53047\ : std_logic;
signal \N__53046\ : std_logic;
signal \N__53045\ : std_logic;
signal \N__53038\ : std_logic;
signal \N__53037\ : std_logic;
signal \N__53036\ : std_logic;
signal \N__53029\ : std_logic;
signal \N__53028\ : std_logic;
signal \N__53027\ : std_logic;
signal \N__53020\ : std_logic;
signal \N__53019\ : std_logic;
signal \N__53018\ : std_logic;
signal \N__53011\ : std_logic;
signal \N__53010\ : std_logic;
signal \N__53009\ : std_logic;
signal \N__53002\ : std_logic;
signal \N__53001\ : std_logic;
signal \N__53000\ : std_logic;
signal \N__52993\ : std_logic;
signal \N__52992\ : std_logic;
signal \N__52991\ : std_logic;
signal \N__52984\ : std_logic;
signal \N__52983\ : std_logic;
signal \N__52982\ : std_logic;
signal \N__52975\ : std_logic;
signal \N__52974\ : std_logic;
signal \N__52973\ : std_logic;
signal \N__52966\ : std_logic;
signal \N__52965\ : std_logic;
signal \N__52964\ : std_logic;
signal \N__52947\ : std_logic;
signal \N__52944\ : std_logic;
signal \N__52941\ : std_logic;
signal \N__52940\ : std_logic;
signal \N__52939\ : std_logic;
signal \N__52936\ : std_logic;
signal \N__52933\ : std_logic;
signal \N__52930\ : std_logic;
signal \N__52929\ : std_logic;
signal \N__52926\ : std_logic;
signal \N__52921\ : std_logic;
signal \N__52918\ : std_logic;
signal \N__52915\ : std_logic;
signal \N__52910\ : std_logic;
signal \N__52905\ : std_logic;
signal \N__52902\ : std_logic;
signal \N__52899\ : std_logic;
signal \N__52896\ : std_logic;
signal \N__52895\ : std_logic;
signal \N__52892\ : std_logic;
signal \N__52889\ : std_logic;
signal \N__52886\ : std_logic;
signal \N__52883\ : std_logic;
signal \N__52878\ : std_logic;
signal \N__52875\ : std_logic;
signal \N__52872\ : std_logic;
signal \N__52869\ : std_logic;
signal \N__52866\ : std_logic;
signal \N__52863\ : std_logic;
signal \N__52862\ : std_logic;
signal \N__52861\ : std_logic;
signal \N__52858\ : std_logic;
signal \N__52853\ : std_logic;
signal \N__52848\ : std_logic;
signal \N__52845\ : std_logic;
signal \N__52842\ : std_logic;
signal \N__52839\ : std_logic;
signal \N__52836\ : std_logic;
signal \N__52833\ : std_logic;
signal \N__52830\ : std_logic;
signal \N__52827\ : std_logic;
signal \N__52826\ : std_logic;
signal \N__52825\ : std_logic;
signal \N__52822\ : std_logic;
signal \N__52819\ : std_logic;
signal \N__52816\ : std_logic;
signal \N__52813\ : std_logic;
signal \N__52810\ : std_logic;
signal \N__52807\ : std_logic;
signal \N__52804\ : std_logic;
signal \N__52799\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52791\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52781\ : std_logic;
signal \N__52778\ : std_logic;
signal \N__52775\ : std_logic;
signal \N__52774\ : std_logic;
signal \N__52771\ : std_logic;
signal \N__52768\ : std_logic;
signal \N__52765\ : std_logic;
signal \N__52762\ : std_logic;
signal \N__52757\ : std_logic;
signal \N__52754\ : std_logic;
signal \N__52751\ : std_logic;
signal \N__52746\ : std_logic;
signal \N__52743\ : std_logic;
signal \N__52740\ : std_logic;
signal \N__52737\ : std_logic;
signal \N__52734\ : std_logic;
signal \N__52731\ : std_logic;
signal \N__52728\ : std_logic;
signal \N__52727\ : std_logic;
signal \N__52726\ : std_logic;
signal \N__52723\ : std_logic;
signal \N__52720\ : std_logic;
signal \N__52717\ : std_logic;
signal \N__52710\ : std_logic;
signal \N__52707\ : std_logic;
signal \N__52704\ : std_logic;
signal \N__52701\ : std_logic;
signal \N__52698\ : std_logic;
signal \N__52695\ : std_logic;
signal \N__52692\ : std_logic;
signal \N__52691\ : std_logic;
signal \N__52690\ : std_logic;
signal \N__52689\ : std_logic;
signal \N__52688\ : std_logic;
signal \N__52687\ : std_logic;
signal \N__52684\ : std_logic;
signal \N__52673\ : std_logic;
signal \N__52672\ : std_logic;
signal \N__52669\ : std_logic;
signal \N__52666\ : std_logic;
signal \N__52663\ : std_logic;
signal \N__52656\ : std_logic;
signal \N__52653\ : std_logic;
signal \N__52650\ : std_logic;
signal \N__52649\ : std_logic;
signal \N__52648\ : std_logic;
signal \N__52647\ : std_logic;
signal \N__52646\ : std_logic;
signal \N__52635\ : std_logic;
signal \N__52634\ : std_logic;
signal \N__52631\ : std_logic;
signal \N__52628\ : std_logic;
signal \N__52627\ : std_logic;
signal \N__52626\ : std_logic;
signal \N__52625\ : std_logic;
signal \N__52624\ : std_logic;
signal \N__52621\ : std_logic;
signal \N__52618\ : std_logic;
signal \N__52609\ : std_logic;
signal \N__52606\ : std_logic;
signal \N__52603\ : std_logic;
signal \N__52600\ : std_logic;
signal \N__52593\ : std_logic;
signal \N__52590\ : std_logic;
signal \N__52589\ : std_logic;
signal \N__52588\ : std_logic;
signal \N__52587\ : std_logic;
signal \N__52586\ : std_logic;
signal \N__52583\ : std_logic;
signal \N__52580\ : std_logic;
signal \N__52577\ : std_logic;
signal \N__52566\ : std_logic;
signal \N__52563\ : std_logic;
signal \N__52562\ : std_logic;
signal \N__52561\ : std_logic;
signal \N__52560\ : std_logic;
signal \N__52557\ : std_logic;
signal \N__52552\ : std_logic;
signal \N__52549\ : std_logic;
signal \N__52542\ : std_logic;
signal \N__52539\ : std_logic;
signal \N__52536\ : std_logic;
signal \N__52533\ : std_logic;
signal \N__52532\ : std_logic;
signal \N__52531\ : std_logic;
signal \N__52528\ : std_logic;
signal \N__52523\ : std_logic;
signal \N__52518\ : std_logic;
signal \N__52515\ : std_logic;
signal \N__52512\ : std_logic;
signal \N__52509\ : std_logic;
signal \N__52506\ : std_logic;
signal \N__52503\ : std_logic;
signal \N__52500\ : std_logic;
signal \N__52499\ : std_logic;
signal \N__52498\ : std_logic;
signal \N__52497\ : std_logic;
signal \N__52496\ : std_logic;
signal \N__52495\ : std_logic;
signal \N__52494\ : std_logic;
signal \N__52493\ : std_logic;
signal \N__52492\ : std_logic;
signal \N__52491\ : std_logic;
signal \N__52490\ : std_logic;
signal \N__52489\ : std_logic;
signal \N__52488\ : std_logic;
signal \N__52487\ : std_logic;
signal \N__52486\ : std_logic;
signal \N__52485\ : std_logic;
signal \N__52484\ : std_logic;
signal \N__52483\ : std_logic;
signal \N__52482\ : std_logic;
signal \N__52481\ : std_logic;
signal \N__52480\ : std_logic;
signal \N__52479\ : std_logic;
signal \N__52478\ : std_logic;
signal \N__52477\ : std_logic;
signal \N__52476\ : std_logic;
signal \N__52475\ : std_logic;
signal \N__52474\ : std_logic;
signal \N__52473\ : std_logic;
signal \N__52472\ : std_logic;
signal \N__52471\ : std_logic;
signal \N__52470\ : std_logic;
signal \N__52469\ : std_logic;
signal \N__52468\ : std_logic;
signal \N__52467\ : std_logic;
signal \N__52466\ : std_logic;
signal \N__52465\ : std_logic;
signal \N__52464\ : std_logic;
signal \N__52463\ : std_logic;
signal \N__52462\ : std_logic;
signal \N__52461\ : std_logic;
signal \N__52460\ : std_logic;
signal \N__52459\ : std_logic;
signal \N__52458\ : std_logic;
signal \N__52457\ : std_logic;
signal \N__52456\ : std_logic;
signal \N__52455\ : std_logic;
signal \N__52454\ : std_logic;
signal \N__52453\ : std_logic;
signal \N__52452\ : std_logic;
signal \N__52451\ : std_logic;
signal \N__52450\ : std_logic;
signal \N__52449\ : std_logic;
signal \N__52448\ : std_logic;
signal \N__52447\ : std_logic;
signal \N__52446\ : std_logic;
signal \N__52445\ : std_logic;
signal \N__52444\ : std_logic;
signal \N__52443\ : std_logic;
signal \N__52442\ : std_logic;
signal \N__52441\ : std_logic;
signal \N__52440\ : std_logic;
signal \N__52439\ : std_logic;
signal \N__52438\ : std_logic;
signal \N__52437\ : std_logic;
signal \N__52436\ : std_logic;
signal \N__52435\ : std_logic;
signal \N__52434\ : std_logic;
signal \N__52433\ : std_logic;
signal \N__52432\ : std_logic;
signal \N__52431\ : std_logic;
signal \N__52430\ : std_logic;
signal \N__52429\ : std_logic;
signal \N__52428\ : std_logic;
signal \N__52427\ : std_logic;
signal \N__52426\ : std_logic;
signal \N__52425\ : std_logic;
signal \N__52424\ : std_logic;
signal \N__52423\ : std_logic;
signal \N__52422\ : std_logic;
signal \N__52421\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52419\ : std_logic;
signal \N__52418\ : std_logic;
signal \N__52417\ : std_logic;
signal \N__52416\ : std_logic;
signal \N__52415\ : std_logic;
signal \N__52414\ : std_logic;
signal \N__52413\ : std_logic;
signal \N__52412\ : std_logic;
signal \N__52411\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52409\ : std_logic;
signal \N__52408\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52406\ : std_logic;
signal \N__52405\ : std_logic;
signal \N__52404\ : std_logic;
signal \N__52403\ : std_logic;
signal \N__52402\ : std_logic;
signal \N__52401\ : std_logic;
signal \N__52400\ : std_logic;
signal \N__52399\ : std_logic;
signal \N__52398\ : std_logic;
signal \N__52397\ : std_logic;
signal \N__52396\ : std_logic;
signal \N__52395\ : std_logic;
signal \N__52394\ : std_logic;
signal \N__52393\ : std_logic;
signal \N__52392\ : std_logic;
signal \N__52391\ : std_logic;
signal \N__52390\ : std_logic;
signal \N__52389\ : std_logic;
signal \N__52388\ : std_logic;
signal \N__52387\ : std_logic;
signal \N__52386\ : std_logic;
signal \N__52385\ : std_logic;
signal \N__52384\ : std_logic;
signal \N__52383\ : std_logic;
signal \N__52382\ : std_logic;
signal \N__52381\ : std_logic;
signal \N__52380\ : std_logic;
signal \N__52379\ : std_logic;
signal \N__52378\ : std_logic;
signal \N__52377\ : std_logic;
signal \N__52376\ : std_logic;
signal \N__52375\ : std_logic;
signal \N__52374\ : std_logic;
signal \N__52373\ : std_logic;
signal \N__52372\ : std_logic;
signal \N__52371\ : std_logic;
signal \N__52370\ : std_logic;
signal \N__52369\ : std_logic;
signal \N__52368\ : std_logic;
signal \N__52367\ : std_logic;
signal \N__52366\ : std_logic;
signal \N__52365\ : std_logic;
signal \N__52092\ : std_logic;
signal \N__52089\ : std_logic;
signal \N__52088\ : std_logic;
signal \N__52087\ : std_logic;
signal \N__52086\ : std_logic;
signal \N__52085\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52083\ : std_logic;
signal \N__52082\ : std_logic;
signal \N__52079\ : std_logic;
signal \N__52076\ : std_logic;
signal \N__52073\ : std_logic;
signal \N__52070\ : std_logic;
signal \N__52067\ : std_logic;
signal \N__52064\ : std_logic;
signal \N__52061\ : std_logic;
signal \N__52058\ : std_logic;
signal \N__52055\ : std_logic;
signal \N__52052\ : std_logic;
signal \N__52049\ : std_logic;
signal \N__52048\ : std_logic;
signal \N__52047\ : std_logic;
signal \N__52046\ : std_logic;
signal \N__52045\ : std_logic;
signal \N__52044\ : std_logic;
signal \N__52043\ : std_logic;
signal \N__52042\ : std_logic;
signal \N__52041\ : std_logic;
signal \N__52040\ : std_logic;
signal \N__52039\ : std_logic;
signal \N__52038\ : std_logic;
signal \N__52037\ : std_logic;
signal \N__52036\ : std_logic;
signal \N__52035\ : std_logic;
signal \N__52034\ : std_logic;
signal \N__52033\ : std_logic;
signal \N__52032\ : std_logic;
signal \N__52031\ : std_logic;
signal \N__52030\ : std_logic;
signal \N__52027\ : std_logic;
signal \N__52026\ : std_logic;
signal \N__52025\ : std_logic;
signal \N__52024\ : std_logic;
signal \N__52023\ : std_logic;
signal \N__52022\ : std_logic;
signal \N__52021\ : std_logic;
signal \N__52020\ : std_logic;
signal \N__52019\ : std_logic;
signal \N__52018\ : std_logic;
signal \N__52017\ : std_logic;
signal \N__52016\ : std_logic;
signal \N__52015\ : std_logic;
signal \N__52014\ : std_logic;
signal \N__52013\ : std_logic;
signal \N__52012\ : std_logic;
signal \N__52011\ : std_logic;
signal \N__52010\ : std_logic;
signal \N__52009\ : std_logic;
signal \N__52008\ : std_logic;
signal \N__52007\ : std_logic;
signal \N__52006\ : std_logic;
signal \N__52005\ : std_logic;
signal \N__52004\ : std_logic;
signal \N__52003\ : std_logic;
signal \N__52002\ : std_logic;
signal \N__52001\ : std_logic;
signal \N__52000\ : std_logic;
signal \N__51999\ : std_logic;
signal \N__51998\ : std_logic;
signal \N__51997\ : std_logic;
signal \N__51996\ : std_logic;
signal \N__51995\ : std_logic;
signal \N__51994\ : std_logic;
signal \N__51993\ : std_logic;
signal \N__51992\ : std_logic;
signal \N__51991\ : std_logic;
signal \N__51990\ : std_logic;
signal \N__51989\ : std_logic;
signal \N__51988\ : std_logic;
signal \N__51987\ : std_logic;
signal \N__51986\ : std_logic;
signal \N__51983\ : std_logic;
signal \N__51982\ : std_logic;
signal \N__51981\ : std_logic;
signal \N__51980\ : std_logic;
signal \N__51979\ : std_logic;
signal \N__51978\ : std_logic;
signal \N__51977\ : std_logic;
signal \N__51976\ : std_logic;
signal \N__51975\ : std_logic;
signal \N__51974\ : std_logic;
signal \N__51973\ : std_logic;
signal \N__51972\ : std_logic;
signal \N__51971\ : std_logic;
signal \N__51970\ : std_logic;
signal \N__51969\ : std_logic;
signal \N__51968\ : std_logic;
signal \N__51967\ : std_logic;
signal \N__51966\ : std_logic;
signal \N__51965\ : std_logic;
signal \N__51964\ : std_logic;
signal \N__51963\ : std_logic;
signal \N__51962\ : std_logic;
signal \N__51961\ : std_logic;
signal \N__51960\ : std_logic;
signal \N__51959\ : std_logic;
signal \N__51958\ : std_logic;
signal \N__51957\ : std_logic;
signal \N__51956\ : std_logic;
signal \N__51955\ : std_logic;
signal \N__51954\ : std_logic;
signal \N__51953\ : std_logic;
signal \N__51952\ : std_logic;
signal \N__51951\ : std_logic;
signal \N__51948\ : std_logic;
signal \N__51947\ : std_logic;
signal \N__51946\ : std_logic;
signal \N__51945\ : std_logic;
signal \N__51944\ : std_logic;
signal \N__51943\ : std_logic;
signal \N__51942\ : std_logic;
signal \N__51941\ : std_logic;
signal \N__51940\ : std_logic;
signal \N__51939\ : std_logic;
signal \N__51936\ : std_logic;
signal \N__51935\ : std_logic;
signal \N__51934\ : std_logic;
signal \N__51933\ : std_logic;
signal \N__51932\ : std_logic;
signal \N__51929\ : std_logic;
signal \N__51928\ : std_logic;
signal \N__51699\ : std_logic;
signal \N__51696\ : std_logic;
signal \N__51693\ : std_logic;
signal \N__51690\ : std_logic;
signal \N__51687\ : std_logic;
signal \N__51684\ : std_logic;
signal \N__51681\ : std_logic;
signal \N__51678\ : std_logic;
signal \N__51677\ : std_logic;
signal \N__51676\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51666\ : std_logic;
signal \N__51663\ : std_logic;
signal \N__51660\ : std_logic;
signal \N__51657\ : std_logic;
signal \N__51654\ : std_logic;
signal \N__51651\ : std_logic;
signal \N__51648\ : std_logic;
signal \N__51645\ : std_logic;
signal \N__51642\ : std_logic;
signal \N__51639\ : std_logic;
signal \N__51636\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51630\ : std_logic;
signal \N__51627\ : std_logic;
signal \N__51624\ : std_logic;
signal \N__51621\ : std_logic;
signal \N__51618\ : std_logic;
signal \N__51615\ : std_logic;
signal \N__51612\ : std_logic;
signal \N__51609\ : std_logic;
signal \N__51606\ : std_logic;
signal \N__51605\ : std_logic;
signal \N__51604\ : std_logic;
signal \N__51597\ : std_logic;
signal \N__51594\ : std_logic;
signal \N__51591\ : std_logic;
signal \N__51588\ : std_logic;
signal \N__51585\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51579\ : std_logic;
signal \N__51576\ : std_logic;
signal \N__51573\ : std_logic;
signal \N__51570\ : std_logic;
signal \N__51567\ : std_logic;
signal \N__51564\ : std_logic;
signal \N__51563\ : std_logic;
signal \N__51562\ : std_logic;
signal \N__51559\ : std_logic;
signal \N__51556\ : std_logic;
signal \N__51553\ : std_logic;
signal \N__51550\ : std_logic;
signal \N__51545\ : std_logic;
signal \N__51542\ : std_logic;
signal \N__51539\ : std_logic;
signal \N__51536\ : std_logic;
signal \N__51533\ : std_logic;
signal \N__51528\ : std_logic;
signal \N__51527\ : std_logic;
signal \N__51524\ : std_logic;
signal \N__51521\ : std_logic;
signal \N__51516\ : std_logic;
signal \N__51513\ : std_logic;
signal \N__51510\ : std_logic;
signal \N__51507\ : std_logic;
signal \N__51504\ : std_logic;
signal \N__51501\ : std_logic;
signal \N__51498\ : std_logic;
signal \N__51497\ : std_logic;
signal \N__51496\ : std_logic;
signal \N__51493\ : std_logic;
signal \N__51490\ : std_logic;
signal \N__51487\ : std_logic;
signal \N__51484\ : std_logic;
signal \N__51481\ : std_logic;
signal \N__51474\ : std_logic;
signal \N__51471\ : std_logic;
signal \N__51468\ : std_logic;
signal \N__51465\ : std_logic;
signal \N__51462\ : std_logic;
signal \N__51459\ : std_logic;
signal \N__51456\ : std_logic;
signal \N__51453\ : std_logic;
signal \N__51450\ : std_logic;
signal \N__51449\ : std_logic;
signal \N__51446\ : std_logic;
signal \N__51443\ : std_logic;
signal \N__51440\ : std_logic;
signal \N__51437\ : std_logic;
signal \N__51434\ : std_logic;
signal \N__51431\ : std_logic;
signal \N__51426\ : std_logic;
signal \N__51425\ : std_logic;
signal \N__51422\ : std_logic;
signal \N__51421\ : std_logic;
signal \N__51418\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51405\ : std_logic;
signal \N__51402\ : std_logic;
signal \N__51399\ : std_logic;
signal \N__51396\ : std_logic;
signal \N__51393\ : std_logic;
signal \N__51390\ : std_logic;
signal \N__51387\ : std_logic;
signal \N__51384\ : std_logic;
signal \N__51381\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51379\ : std_logic;
signal \N__51378\ : std_logic;
signal \N__51375\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51370\ : std_logic;
signal \N__51369\ : std_logic;
signal \N__51368\ : std_logic;
signal \N__51367\ : std_logic;
signal \N__51364\ : std_logic;
signal \N__51361\ : std_logic;
signal \N__51360\ : std_logic;
signal \N__51359\ : std_logic;
signal \N__51358\ : std_logic;
signal \N__51355\ : std_logic;
signal \N__51352\ : std_logic;
signal \N__51349\ : std_logic;
signal \N__51346\ : std_logic;
signal \N__51337\ : std_logic;
signal \N__51328\ : std_logic;
signal \N__51323\ : std_logic;
signal \N__51320\ : std_logic;
signal \N__51317\ : std_logic;
signal \N__51314\ : std_logic;
signal \N__51309\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51299\ : std_logic;
signal \N__51296\ : std_logic;
signal \N__51293\ : std_logic;
signal \N__51290\ : std_logic;
signal \N__51287\ : std_logic;
signal \N__51284\ : std_logic;
signal \N__51279\ : std_logic;
signal \N__51276\ : std_logic;
signal \N__51273\ : std_logic;
signal \N__51270\ : std_logic;
signal \N__51267\ : std_logic;
signal \N__51264\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51260\ : std_logic;
signal \N__51257\ : std_logic;
signal \N__51254\ : std_logic;
signal \N__51253\ : std_logic;
signal \N__51250\ : std_logic;
signal \N__51247\ : std_logic;
signal \N__51244\ : std_logic;
signal \N__51239\ : std_logic;
signal \N__51234\ : std_logic;
signal \N__51231\ : std_logic;
signal \N__51228\ : std_logic;
signal \N__51225\ : std_logic;
signal \N__51222\ : std_logic;
signal \N__51221\ : std_logic;
signal \N__51218\ : std_logic;
signal \N__51215\ : std_logic;
signal \N__51212\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51201\ : std_logic;
signal \N__51198\ : std_logic;
signal \N__51195\ : std_logic;
signal \N__51192\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51190\ : std_logic;
signal \N__51187\ : std_logic;
signal \N__51184\ : std_logic;
signal \N__51181\ : std_logic;
signal \N__51178\ : std_logic;
signal \N__51171\ : std_logic;
signal \N__51168\ : std_logic;
signal \N__51165\ : std_logic;
signal \N__51162\ : std_logic;
signal \N__51159\ : std_logic;
signal \N__51156\ : std_logic;
signal \N__51153\ : std_logic;
signal \N__51150\ : std_logic;
signal \N__51149\ : std_logic;
signal \N__51148\ : std_logic;
signal \N__51145\ : std_logic;
signal \N__51142\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51129\ : std_logic;
signal \N__51126\ : std_logic;
signal \N__51123\ : std_logic;
signal \N__51120\ : std_logic;
signal \N__51117\ : std_logic;
signal \N__51116\ : std_logic;
signal \N__51115\ : std_logic;
signal \N__51112\ : std_logic;
signal \N__51109\ : std_logic;
signal \N__51106\ : std_logic;
signal \N__51103\ : std_logic;
signal \N__51100\ : std_logic;
signal \N__51093\ : std_logic;
signal \N__51090\ : std_logic;
signal \N__51087\ : std_logic;
signal \N__51084\ : std_logic;
signal \N__51081\ : std_logic;
signal \N__51080\ : std_logic;
signal \N__51077\ : std_logic;
signal \N__51074\ : std_logic;
signal \N__51071\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51063\ : std_logic;
signal \N__51060\ : std_logic;
signal \N__51057\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51051\ : std_logic;
signal \N__51048\ : std_logic;
signal \N__51045\ : std_logic;
signal \N__51042\ : std_logic;
signal \N__51039\ : std_logic;
signal \N__51036\ : std_logic;
signal \N__51033\ : std_logic;
signal \N__51030\ : std_logic;
signal \N__51027\ : std_logic;
signal \N__51024\ : std_logic;
signal \N__51021\ : std_logic;
signal \N__51018\ : std_logic;
signal \N__51015\ : std_logic;
signal \N__51012\ : std_logic;
signal \N__51009\ : std_logic;
signal \N__51006\ : std_logic;
signal \N__51003\ : std_logic;
signal \N__51000\ : std_logic;
signal \N__50997\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50991\ : std_logic;
signal \N__50988\ : std_logic;
signal \N__50985\ : std_logic;
signal \N__50982\ : std_logic;
signal \N__50979\ : std_logic;
signal \N__50976\ : std_logic;
signal \N__50973\ : std_logic;
signal \N__50970\ : std_logic;
signal \N__50967\ : std_logic;
signal \N__50964\ : std_logic;
signal \N__50961\ : std_logic;
signal \N__50958\ : std_logic;
signal \N__50955\ : std_logic;
signal \N__50952\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50946\ : std_logic;
signal \N__50943\ : std_logic;
signal \N__50940\ : std_logic;
signal \N__50937\ : std_logic;
signal \N__50934\ : std_logic;
signal \N__50931\ : std_logic;
signal \N__50928\ : std_logic;
signal \N__50925\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50919\ : std_logic;
signal \N__50916\ : std_logic;
signal \N__50913\ : std_logic;
signal \N__50910\ : std_logic;
signal \N__50907\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50901\ : std_logic;
signal \N__50898\ : std_logic;
signal \N__50895\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50891\ : std_logic;
signal \N__50888\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50880\ : std_logic;
signal \N__50879\ : std_logic;
signal \N__50878\ : std_logic;
signal \N__50877\ : std_logic;
signal \N__50876\ : std_logic;
signal \N__50875\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50873\ : std_logic;
signal \N__50870\ : std_logic;
signal \N__50869\ : std_logic;
signal \N__50866\ : std_logic;
signal \N__50861\ : std_logic;
signal \N__50856\ : std_logic;
signal \N__50853\ : std_logic;
signal \N__50852\ : std_logic;
signal \N__50851\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50849\ : std_logic;
signal \N__50848\ : std_logic;
signal \N__50847\ : std_logic;
signal \N__50846\ : std_logic;
signal \N__50845\ : std_logic;
signal \N__50838\ : std_logic;
signal \N__50837\ : std_logic;
signal \N__50836\ : std_logic;
signal \N__50835\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50833\ : std_logic;
signal \N__50826\ : std_logic;
signal \N__50825\ : std_logic;
signal \N__50824\ : std_logic;
signal \N__50823\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50819\ : std_logic;
signal \N__50818\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50816\ : std_logic;
signal \N__50815\ : std_logic;
signal \N__50804\ : std_logic;
signal \N__50799\ : std_logic;
signal \N__50796\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50788\ : std_logic;
signal \N__50785\ : std_logic;
signal \N__50780\ : std_logic;
signal \N__50777\ : std_logic;
signal \N__50768\ : std_logic;
signal \N__50765\ : std_logic;
signal \N__50756\ : std_logic;
signal \N__50751\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50721\ : std_logic;
signal \N__50718\ : std_logic;
signal \N__50715\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50709\ : std_logic;
signal \N__50708\ : std_logic;
signal \N__50705\ : std_logic;
signal \N__50702\ : std_logic;
signal \N__50697\ : std_logic;
signal \N__50696\ : std_logic;
signal \N__50693\ : std_logic;
signal \N__50690\ : std_logic;
signal \N__50687\ : std_logic;
signal \N__50684\ : std_logic;
signal \N__50679\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50672\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50663\ : std_logic;
signal \N__50662\ : std_logic;
signal \N__50657\ : std_logic;
signal \N__50654\ : std_logic;
signal \N__50651\ : std_logic;
signal \N__50646\ : std_logic;
signal \N__50643\ : std_logic;
signal \N__50640\ : std_logic;
signal \N__50639\ : std_logic;
signal \N__50636\ : std_logic;
signal \N__50633\ : std_logic;
signal \N__50628\ : std_logic;
signal \N__50627\ : std_logic;
signal \N__50624\ : std_logic;
signal \N__50621\ : std_logic;
signal \N__50618\ : std_logic;
signal \N__50617\ : std_logic;
signal \N__50612\ : std_logic;
signal \N__50609\ : std_logic;
signal \N__50606\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50598\ : std_logic;
signal \N__50595\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50591\ : std_logic;
signal \N__50588\ : std_logic;
signal \N__50583\ : std_logic;
signal \N__50582\ : std_logic;
signal \N__50579\ : std_logic;
signal \N__50576\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50574\ : std_logic;
signal \N__50573\ : std_logic;
signal \N__50570\ : std_logic;
signal \N__50567\ : std_logic;
signal \N__50564\ : std_logic;
signal \N__50561\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50529\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50511\ : std_logic;
signal \N__50508\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50471\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50460\ : std_logic;
signal \N__50457\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50451\ : std_logic;
signal \N__50448\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50444\ : std_logic;
signal \N__50441\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50433\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50426\ : std_logic;
signal \N__50423\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50415\ : std_logic;
signal \N__50414\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50397\ : std_logic;
signal \N__50396\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50382\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50373\ : std_logic;
signal \N__50370\ : std_logic;
signal \N__50369\ : std_logic;
signal \N__50366\ : std_logic;
signal \N__50363\ : std_logic;
signal \N__50358\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50300\ : std_logic;
signal \N__50297\ : std_logic;
signal \N__50294\ : std_logic;
signal \N__50289\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50273\ : std_logic;
signal \N__50270\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50246\ : std_logic;
signal \N__50243\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50235\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50229\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50225\ : std_logic;
signal \N__50222\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50213\ : std_logic;
signal \N__50208\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50204\ : std_logic;
signal \N__50201\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50193\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50187\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50180\ : std_logic;
signal \N__50177\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50171\ : std_logic;
signal \N__50168\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50156\ : std_logic;
signal \N__50155\ : std_logic;
signal \N__50152\ : std_logic;
signal \N__50149\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50147\ : std_logic;
signal \N__50146\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50141\ : std_logic;
signal \N__50140\ : std_logic;
signal \N__50135\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50125\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50119\ : std_logic;
signal \N__50116\ : std_logic;
signal \N__50113\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50098\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50085\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50071\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50061\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50057\ : std_logic;
signal \N__50054\ : std_logic;
signal \N__50051\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50045\ : std_logic;
signal \N__50040\ : std_logic;
signal \N__50037\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50025\ : std_logic;
signal \N__50022\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50015\ : std_logic;
signal \N__50012\ : std_logic;
signal \N__50009\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49995\ : std_logic;
signal \N__49992\ : std_logic;
signal \N__49991\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49983\ : std_logic;
signal \N__49982\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49976\ : std_logic;
signal \N__49973\ : std_logic;
signal \N__49970\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49961\ : std_logic;
signal \N__49958\ : std_logic;
signal \N__49957\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49938\ : std_logic;
signal \N__49935\ : std_logic;
signal \N__49932\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49926\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49917\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49913\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49904\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49880\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49862\ : std_logic;
signal \N__49859\ : std_logic;
signal \N__49856\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49843\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49826\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49809\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49772\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49766\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49760\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49731\ : std_logic;
signal \N__49728\ : std_logic;
signal \N__49725\ : std_logic;
signal \N__49722\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49716\ : std_logic;
signal \N__49713\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49689\ : std_logic;
signal \N__49686\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49680\ : std_logic;
signal \N__49677\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49668\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49664\ : std_logic;
signal \N__49661\ : std_logic;
signal \N__49658\ : std_logic;
signal \N__49653\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49647\ : std_logic;
signal \N__49644\ : std_logic;
signal \N__49641\ : std_logic;
signal \N__49640\ : std_logic;
signal \N__49637\ : std_logic;
signal \N__49634\ : std_logic;
signal \N__49631\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49617\ : std_logic;
signal \N__49614\ : std_logic;
signal \N__49611\ : std_logic;
signal \N__49610\ : std_logic;
signal \N__49607\ : std_logic;
signal \N__49604\ : std_logic;
signal \N__49599\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49578\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49571\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49557\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49479\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49452\ : std_logic;
signal \N__49449\ : std_logic;
signal \N__49446\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49440\ : std_logic;
signal \N__49437\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49422\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49398\ : std_logic;
signal \N__49395\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49386\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49382\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49355\ : std_logic;
signal \N__49352\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49345\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49335\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49329\ : std_logic;
signal \N__49328\ : std_logic;
signal \N__49325\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49315\ : std_logic;
signal \N__49308\ : std_logic;
signal \N__49305\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49301\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49294\ : std_logic;
signal \N__49291\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49278\ : std_logic;
signal \N__49275\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49271\ : std_logic;
signal \N__49270\ : std_logic;
signal \N__49267\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49261\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49251\ : std_logic;
signal \N__49248\ : std_logic;
signal \N__49247\ : std_logic;
signal \N__49244\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49240\ : std_logic;
signal \N__49237\ : std_logic;
signal \N__49234\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49220\ : std_logic;
signal \N__49219\ : std_logic;
signal \N__49216\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49210\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49196\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49166\ : std_logic;
signal \N__49165\ : std_logic;
signal \N__49162\ : std_logic;
signal \N__49159\ : std_logic;
signal \N__49156\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49097\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49086\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49082\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49070\ : std_logic;
signal \N__49065\ : std_logic;
signal \N__49062\ : std_logic;
signal \N__49059\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49052\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49038\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49036\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49032\ : std_logic;
signal \N__49031\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49029\ : std_logic;
signal \N__49028\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49025\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49022\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49019\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49016\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48971\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48944\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48921\ : std_logic;
signal \N__48918\ : std_logic;
signal \N__48917\ : std_logic;
signal \N__48914\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48908\ : std_logic;
signal \N__48903\ : std_logic;
signal \N__48902\ : std_logic;
signal \N__48899\ : std_logic;
signal \N__48898\ : std_logic;
signal \N__48895\ : std_logic;
signal \N__48892\ : std_logic;
signal \N__48889\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48882\ : std_logic;
signal \N__48879\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48850\ : std_logic;
signal \N__48847\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48828\ : std_logic;
signal \N__48827\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48823\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48807\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48794\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48788\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48761\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48740\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48732\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48725\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48698\ : std_logic;
signal \N__48695\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48675\ : std_logic;
signal \N__48674\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48665\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48657\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48630\ : std_logic;
signal \N__48627\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48603\ : std_logic;
signal \N__48600\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48593\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48560\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48552\ : std_logic;
signal \N__48549\ : std_logic;
signal \N__48546\ : std_logic;
signal \N__48543\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48506\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48485\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48476\ : std_logic;
signal \N__48473\ : std_logic;
signal \N__48470\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48455\ : std_logic;
signal \N__48452\ : std_logic;
signal \N__48449\ : std_logic;
signal \N__48446\ : std_logic;
signal \N__48441\ : std_logic;
signal \N__48438\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48434\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48371\ : std_logic;
signal \N__48368\ : std_logic;
signal \N__48365\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48357\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48353\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48347\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48320\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48309\ : std_logic;
signal \N__48306\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48230\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48114\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48104\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48077\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48053\ : std_logic;
signal \N__48050\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48015\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48008\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47979\ : std_logic;
signal \N__47976\ : std_logic;
signal \N__47975\ : std_logic;
signal \N__47972\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47748\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47667\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47639\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47580\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47574\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47562\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47550\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47529\ : std_logic;
signal \N__47526\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47504\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47262\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47223\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47207\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47187\ : std_logic;
signal \N__47184\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47177\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47043\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46838\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46771\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46721\ : std_logic;
signal \N__46718\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46705\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46685\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46592\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46577\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46548\ : std_logic;
signal \N__46545\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46489\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46486\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46436\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46365\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46357\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46286\ : std_logic;
signal \N__46283\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46187\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46144\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46088\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46073\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45921\ : std_logic;
signal \N__45918\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45855\ : std_logic;
signal \N__45852\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45792\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45764\ : std_logic;
signal \N__45761\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45666\ : std_logic;
signal \N__45663\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45474\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45420\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45395\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45351\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45342\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45237\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45192\ : std_logic;
signal \N__45189\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45171\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44996\ : std_logic;
signal \N__44993\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44814\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44673\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44541\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44511\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44501\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44246\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44192\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44110\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44107\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44104\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44101\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44051\ : std_logic;
signal \N__44048\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44030\ : std_logic;
signal \N__44023\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44002\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43961\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43692\ : std_logic;
signal \N__43689\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43659\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43551\ : std_logic;
signal \N__43548\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43503\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43383\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43374\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43326\ : std_logic;
signal \N__43323\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43197\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43191\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43061\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42935\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42912\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42662\ : std_logic;
signal \N__42659\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42497\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42410\ : std_logic;
signal \N__42407\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42157\ : std_logic;
signal \N__42154\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41930\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41835\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41759\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41590\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41411\ : std_logic;
signal \N__41408\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41352\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41300\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41267\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40816\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40727\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40339\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40295\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39956\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39672\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39299\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39194\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37572\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\ : std_logic;
signal \N_94_i_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_25\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal un8_start_stop : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \bfn_3_11_0_\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \bfn_3_12_0_\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.control_input_cry_13\ : std_logic;
signal \current_shift_inst.control_input_cry_14\ : std_logic;
signal \current_shift_inst.control_input_cry_15\ : std_logic;
signal \bfn_3_13_0_\ : std_logic;
signal \current_shift_inst.control_input_cry_16\ : std_logic;
signal \current_shift_inst.control_input_cry_17\ : std_logic;
signal \current_shift_inst.control_input_cry_18\ : std_logic;
signal \current_shift_inst.control_input_cry_19\ : std_logic;
signal \current_shift_inst.control_input_cry_20\ : std_logic;
signal \current_shift_inst.control_input_cry_21\ : std_logic;
signal \current_shift_inst.control_input_cry_22\ : std_logic;
signal \current_shift_inst.control_input_cry_23\ : std_logic;
signal \bfn_3_14_0_\ : std_logic;
signal \current_shift_inst.control_input_cry_24\ : std_logic;
signal \current_shift_inst.control_input_cry_25\ : std_logic;
signal \current_shift_inst.control_input_cry_26\ : std_logic;
signal \current_shift_inst.control_input_cry_27\ : std_logic;
signal \current_shift_inst.control_input_cry_28\ : std_logic;
signal \current_shift_inst.control_input_cry_29\ : std_logic;
signal \current_shift_inst.control_input_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44_cascade_\ : std_logic;
signal \current_shift_inst.N_1571_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_77\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \current_shift_inst.control_input_axb_13\ : std_logic;
signal \current_shift_inst.control_input_axb_18\ : std_logic;
signal \current_shift_inst.control_input_axb_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.control_input_axb_27\ : std_logic;
signal \current_shift_inst.control_input_axb_22\ : std_logic;
signal \current_shift_inst.control_input_axb_24\ : std_logic;
signal \current_shift_inst.control_input_axb_23\ : std_logic;
signal \current_shift_inst.control_input_axb_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.control_input_axb_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_16_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.control_input_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_29\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_30\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.control_input_axb_14\ : std_logic;
signal \current_shift_inst.control_input_axb_26\ : std_logic;
signal \current_shift_inst.control_input_axb_21\ : std_logic;
signal \current_shift_inst.control_input_axb_17\ : std_logic;
signal \current_shift_inst.control_input_axb_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_22\ : std_logic;
signal \current_shift_inst.control_input_axb_16\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.control_input_axb_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_28\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst2.start_flagZ0\ : std_logic;
signal \phase_controller_inst2.state_ns_0_0_1\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_8\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_16\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_axb_28\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_8\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_16\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_19\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_8_22_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal s4_phy_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_start_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal s3_phy_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_0_sqmuxa\ : std_logic;
signal \bfn_10_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_7\ : std_logic;
signal \bfn_10_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_15\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_23\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_i_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0_g\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_10_20_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_start_0\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_0\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_8\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_15\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_30\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \bfn_11_21_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_0\ : std_logic;
signal \bfn_11_25_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_8\ : std_logic;
signal \bfn_11_26_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_15\ : std_logic;
signal \bfn_11_27_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_30\ : std_logic;
signal \bfn_11_28_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt24\ : std_logic;
signal \current_shift_inst.timer_s1.N_154_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt26\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_14\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.timer_s1.N_153_i_g\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ1Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_0\ : std_logic;
signal \bfn_12_27_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_8\ : std_logic;
signal \bfn_12_28_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_15\ : std_logic;
signal \bfn_12_29_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_24\ : std_logic;
signal \bfn_12_30_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_i_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0_g\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_7\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_15\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_23\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_i_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal il_max_comp1_c : std_logic;
signal start_stop_c : std_logic;
signal \phase_controller_inst1.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst1.state_ns_0_0_1_cascade_\ : std_logic;
signal \phase_controller_inst1.start_flagZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_start_0\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.measured_delay_tr_i_31\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_1 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_2 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_3 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_4 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_5 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_6 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_7 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_8 : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_9 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_10 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_11 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_12 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_13 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_14 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_15 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_16 : std_logic;
signal \bfn_13_21_0_\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_17 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_18 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_20 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_21 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_22 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_23 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_24 : std_logic;
signal \bfn_13_22_0_\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_25 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_26 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_27 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_13_25_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_13_26_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_158_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_19 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt18\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \current_shift_inst.timer_s1.N_153_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_0\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_8\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_15\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_30\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_0\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_8\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_15\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_30\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_0\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_8\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_15\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_23\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_i_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0\ : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_28 : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_14_25_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_14_26_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_14_27_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal s1_phy_c : std_logic;
signal state_3 : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ1Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \elapsed_time_ns_1_RNIDC91B_0_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_157_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \elapsed_time_ns_1_RNIED91B_0_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\ : std_logic;
signal \bfn_15_28_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \bfn_15_29_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \bfn_15_30_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_16_24_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_15\ : std_logic;
signal pwm_duty_input_10 : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_4\ : std_logic;
signal \bfn_16_28_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_23\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\ : std_logic;
signal \bfn_16_29_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_16_30_0_\ : std_logic;
signal \GB_BUFFER_red_c_g_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.measured_delay_hc_i_31\ : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_1 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_2 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_3 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_4 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_5 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_6 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_7 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_8 : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_9 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_10 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_11 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_12 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_13 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_14 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_15 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_20 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_21 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_22 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_23 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27\ : std_logic;
signal \elapsed_time_ns_1_RNIDV2T9_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \elapsed_time_ns_1_RNIE03T9_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_28 : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_17_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_17_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_17_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_156_i\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_17_24_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_17_25_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \pwm_generator_inst.un19_threshold_0_axb_0\ : std_logic;
signal \pwm_generator_inst.un14_counter_0\ : std_logic;
signal \bfn_17_26_0_\ : std_logic;
signal \pwm_generator_inst.un14_counter_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_axb_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_axb_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_cry_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_axb_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_cry_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_axb_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_cry_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_8\ : std_logic;
signal \bfn_17_27_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_axb_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_axb_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_axb_8\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_16 : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_18 : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_19 : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_17 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_27 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_27\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_26 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_26\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_24 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_24\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_25 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_155_i\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_0\ : std_logic;
signal \bfn_20_25_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_8\ : std_logic;
signal \bfn_20_26_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \pwm_generator_inst.un19_threshold_0_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_20_27_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal \current_shift_inst.PI_CTRL.N_152\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal pwm_duty_input_1 : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_94\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal pwm_duty_input_8 : std_logic;
signal \current_shift_inst.PI_CTRL.N_150\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal pwm_output_wire : std_logic;
signal s2_phy_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    pwm_output <= pwm_output_wire;
    s2_phy <= s2_phy_wire;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    il_max_comp1_wire <= il_max_comp1;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ <= \N__23358\&\N__23235\&\N__23990\&\N__23211\&\N__23406\&\N__23187\&\N__23439\&\N__23807\&\N__23723\&\N__23837\&\N__23490\&\N__23259\&\N__23463\&\N__23379\&\N__23064\&\N__26103\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__46144\&'0'&\N__46143\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__44966\&\N__44959\&\N__44964\&\N__44958\&\N__44965\&\N__44957\&\N__44967\&\N__44954\&\N__44960\&\N__44953\&\N__44961\&\N__44955\&\N__44962\&\N__44956\&\N__44963\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__46448\&\N__46445\&'0'&'0'&'0'&\N__46443\&\N__46447\&\N__46444\&\N__46446\;
    \pwm_generator_inst.un2_threshold_2_1_16\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_2_1_15\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_2_14\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_2_13\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ <= '0'&\N__44968\&\N__44971\&\N__44969\&\N__44972\&\N__44970\&\N__52836\&\N__52701\&\N__52509\&\N__52791\&\N__52743\&\N__52878\&\N__51510\&\N__51633\&\N__51576\&\N__51615\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__46585\&\N__46582\&'0'&'0'&'0'&\N__46580\&\N__46584\&\N__46581\&\N__46583\;
    \pwm_generator_inst.un2_threshold_1_25\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_1_24\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_1_23\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_1_22\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_1_21\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_1_20\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(0);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ <= '0'&\N__23280\&\N__26082\&\N__23297\&\N__26117\&\N__23319\&\N__23855\&\N__23882\&\N__23088\&\N__23622\&\N__26150\&\N__23777\&\N__23517\&\N__23915\&\N__23741\&\N__22673\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__46307\&'0'&\N__46306\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(19);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(18);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(17);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(16);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.un1_integrator\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__21981\,
            RESETB => \N__45795\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__46145\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__46142\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__46449\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__46442\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__46586\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__46579\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__46305\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__46304\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__53074\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53076\,
            DIN => \N__53075\,
            DOUT => \N__53074\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53076\,
            PADOUT => \N__53075\,
            PADIN => \N__53074\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53065\,
            DIN => \N__53064\,
            DOUT => \N__53063\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53065\,
            PADOUT => \N__53064\,
            PADIN => \N__53063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__49554\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53056\,
            DIN => \N__53055\,
            DOUT => \N__53054\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53056\,
            PADOUT => \N__53055\,
            PADIN => \N__53054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__38235\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53047\,
            DIN => \N__53046\,
            DOUT => \N__53045\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53047\,
            PADOUT => \N__53046\,
            PADIN => \N__53045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53038\,
            DIN => \N__53037\,
            DOUT => \N__53036\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53038\,
            PADOUT => \N__53037\,
            PADIN => \N__53036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__41250\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53029\,
            DIN => \N__53028\,
            DOUT => \N__53027\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53029\,
            PADOUT => \N__53028\,
            PADIN => \N__53027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25044\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53020\,
            DIN => \N__53019\,
            DOUT => \N__53018\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53020\,
            PADOUT => \N__53019\,
            PADIN => \N__53018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53011\,
            DIN => \N__53010\,
            DOUT => \N__53009\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53011\,
            PADOUT => \N__53010\,
            PADIN => \N__53009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25812\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53002\,
            DIN => \N__53001\,
            DOUT => \N__53000\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53002\,
            PADOUT => \N__53001\,
            PADIN => \N__53000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52993\,
            DIN => \N__52992\,
            DOUT => \N__52991\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52993\,
            PADOUT => \N__52992\,
            PADIN => \N__52991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52984\,
            DIN => \N__52983\,
            DOUT => \N__52982\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52984\,
            PADOUT => \N__52983\,
            PADIN => \N__52982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52975\,
            DIN => \N__52974\,
            DOUT => \N__52973\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52975\,
            PADOUT => \N__52974\,
            PADIN => \N__52973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52966\,
            DIN => \N__52965\,
            DOUT => \N__52964\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52966\,
            PADOUT => \N__52965\,
            PADIN => \N__52964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__12380\ : InMux
    port map (
            O => \N__52947\,
            I => \N__52944\
        );

    \I__12379\ : LocalMux
    port map (
            O => \N__52944\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__12378\ : InMux
    port map (
            O => \N__52941\,
            I => \N__52936\
        );

    \I__12377\ : CascadeMux
    port map (
            O => \N__52940\,
            I => \N__52933\
        );

    \I__12376\ : CascadeMux
    port map (
            O => \N__52939\,
            I => \N__52930\
        );

    \I__12375\ : LocalMux
    port map (
            O => \N__52936\,
            I => \N__52926\
        );

    \I__12374\ : InMux
    port map (
            O => \N__52933\,
            I => \N__52921\
        );

    \I__12373\ : InMux
    port map (
            O => \N__52930\,
            I => \N__52921\
        );

    \I__12372\ : InMux
    port map (
            O => \N__52929\,
            I => \N__52918\
        );

    \I__12371\ : Span4Mux_v
    port map (
            O => \N__52926\,
            I => \N__52915\
        );

    \I__12370\ : LocalMux
    port map (
            O => \N__52921\,
            I => \N__52910\
        );

    \I__12369\ : LocalMux
    port map (
            O => \N__52918\,
            I => \N__52910\
        );

    \I__12368\ : Sp12to4
    port map (
            O => \N__52915\,
            I => \N__52905\
        );

    \I__12367\ : Span12Mux_v
    port map (
            O => \N__52910\,
            I => \N__52905\
        );

    \I__12366\ : Span12Mux_h
    port map (
            O => \N__52905\,
            I => \N__52902\
        );

    \I__12365\ : Odrv12
    port map (
            O => \N__52902\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__12364\ : CascadeMux
    port map (
            O => \N__52899\,
            I => \N__52896\
        );

    \I__12363\ : InMux
    port map (
            O => \N__52896\,
            I => \N__52892\
        );

    \I__12362\ : CascadeMux
    port map (
            O => \N__52895\,
            I => \N__52889\
        );

    \I__12361\ : LocalMux
    port map (
            O => \N__52892\,
            I => \N__52886\
        );

    \I__12360\ : InMux
    port map (
            O => \N__52889\,
            I => \N__52883\
        );

    \I__12359\ : Odrv4
    port map (
            O => \N__52886\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__12358\ : LocalMux
    port map (
            O => \N__52883\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__12357\ : InMux
    port map (
            O => \N__52878\,
            I => \N__52875\
        );

    \I__12356\ : LocalMux
    port map (
            O => \N__52875\,
            I => \N__52872\
        );

    \I__12355\ : Odrv4
    port map (
            O => \N__52872\,
            I => pwm_duty_input_4
        );

    \I__12354\ : CascadeMux
    port map (
            O => \N__52869\,
            I => \N__52866\
        );

    \I__12353\ : InMux
    port map (
            O => \N__52866\,
            I => \N__52863\
        );

    \I__12352\ : LocalMux
    port map (
            O => \N__52863\,
            I => \N__52858\
        );

    \I__12351\ : InMux
    port map (
            O => \N__52862\,
            I => \N__52853\
        );

    \I__12350\ : InMux
    port map (
            O => \N__52861\,
            I => \N__52853\
        );

    \I__12349\ : Span4Mux_v
    port map (
            O => \N__52858\,
            I => \N__52848\
        );

    \I__12348\ : LocalMux
    port map (
            O => \N__52853\,
            I => \N__52848\
        );

    \I__12347\ : Span4Mux_h
    port map (
            O => \N__52848\,
            I => \N__52845\
        );

    \I__12346\ : Span4Mux_h
    port map (
            O => \N__52845\,
            I => \N__52842\
        );

    \I__12345\ : Span4Mux_h
    port map (
            O => \N__52842\,
            I => \N__52839\
        );

    \I__12344\ : Odrv4
    port map (
            O => \N__52839\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__12343\ : InMux
    port map (
            O => \N__52836\,
            I => \N__52833\
        );

    \I__12342\ : LocalMux
    port map (
            O => \N__52833\,
            I => \N__52830\
        );

    \I__12341\ : Odrv4
    port map (
            O => \N__52830\,
            I => pwm_duty_input_9
        );

    \I__12340\ : InMux
    port map (
            O => \N__52827\,
            I => \N__52822\
        );

    \I__12339\ : CascadeMux
    port map (
            O => \N__52826\,
            I => \N__52819\
        );

    \I__12338\ : InMux
    port map (
            O => \N__52825\,
            I => \N__52816\
        );

    \I__12337\ : LocalMux
    port map (
            O => \N__52822\,
            I => \N__52813\
        );

    \I__12336\ : InMux
    port map (
            O => \N__52819\,
            I => \N__52810\
        );

    \I__12335\ : LocalMux
    port map (
            O => \N__52816\,
            I => \N__52807\
        );

    \I__12334\ : Span4Mux_v
    port map (
            O => \N__52813\,
            I => \N__52804\
        );

    \I__12333\ : LocalMux
    port map (
            O => \N__52810\,
            I => \N__52799\
        );

    \I__12332\ : Sp12to4
    port map (
            O => \N__52807\,
            I => \N__52799\
        );

    \I__12331\ : Sp12to4
    port map (
            O => \N__52804\,
            I => \N__52794\
        );

    \I__12330\ : Span12Mux_s11_v
    port map (
            O => \N__52799\,
            I => \N__52794\
        );

    \I__12329\ : Odrv12
    port map (
            O => \N__52794\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__12328\ : InMux
    port map (
            O => \N__52791\,
            I => \N__52788\
        );

    \I__12327\ : LocalMux
    port map (
            O => \N__52788\,
            I => \N__52785\
        );

    \I__12326\ : Odrv4
    port map (
            O => \N__52785\,
            I => pwm_duty_input_6
        );

    \I__12325\ : CascadeMux
    port map (
            O => \N__52782\,
            I => \N__52778\
        );

    \I__12324\ : CascadeMux
    port map (
            O => \N__52781\,
            I => \N__52775\
        );

    \I__12323\ : InMux
    port map (
            O => \N__52778\,
            I => \N__52771\
        );

    \I__12322\ : InMux
    port map (
            O => \N__52775\,
            I => \N__52768\
        );

    \I__12321\ : InMux
    port map (
            O => \N__52774\,
            I => \N__52765\
        );

    \I__12320\ : LocalMux
    port map (
            O => \N__52771\,
            I => \N__52762\
        );

    \I__12319\ : LocalMux
    port map (
            O => \N__52768\,
            I => \N__52757\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__52765\,
            I => \N__52757\
        );

    \I__12317\ : Span4Mux_v
    port map (
            O => \N__52762\,
            I => \N__52754\
        );

    \I__12316\ : Span4Mux_v
    port map (
            O => \N__52757\,
            I => \N__52751\
        );

    \I__12315\ : Sp12to4
    port map (
            O => \N__52754\,
            I => \N__52746\
        );

    \I__12314\ : Sp12to4
    port map (
            O => \N__52751\,
            I => \N__52746\
        );

    \I__12313\ : Odrv12
    port map (
            O => \N__52746\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__12312\ : InMux
    port map (
            O => \N__52743\,
            I => \N__52740\
        );

    \I__12311\ : LocalMux
    port map (
            O => \N__52740\,
            I => \N__52737\
        );

    \I__12310\ : Span4Mux_v
    port map (
            O => \N__52737\,
            I => \N__52734\
        );

    \I__12309\ : Odrv4
    port map (
            O => \N__52734\,
            I => pwm_duty_input_5
        );

    \I__12308\ : InMux
    port map (
            O => \N__52731\,
            I => \N__52728\
        );

    \I__12307\ : LocalMux
    port map (
            O => \N__52728\,
            I => \N__52723\
        );

    \I__12306\ : InMux
    port map (
            O => \N__52727\,
            I => \N__52720\
        );

    \I__12305\ : InMux
    port map (
            O => \N__52726\,
            I => \N__52717\
        );

    \I__12304\ : Span4Mux_s3_h
    port map (
            O => \N__52723\,
            I => \N__52710\
        );

    \I__12303\ : LocalMux
    port map (
            O => \N__52720\,
            I => \N__52710\
        );

    \I__12302\ : LocalMux
    port map (
            O => \N__52717\,
            I => \N__52710\
        );

    \I__12301\ : Span4Mux_v
    port map (
            O => \N__52710\,
            I => \N__52707\
        );

    \I__12300\ : Sp12to4
    port map (
            O => \N__52707\,
            I => \N__52704\
        );

    \I__12299\ : Odrv12
    port map (
            O => \N__52704\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__12298\ : InMux
    port map (
            O => \N__52701\,
            I => \N__52698\
        );

    \I__12297\ : LocalMux
    port map (
            O => \N__52698\,
            I => \N__52695\
        );

    \I__12296\ : Odrv4
    port map (
            O => \N__52695\,
            I => pwm_duty_input_8
        );

    \I__12295\ : InMux
    port map (
            O => \N__52692\,
            I => \N__52684\
        );

    \I__12294\ : InMux
    port map (
            O => \N__52691\,
            I => \N__52673\
        );

    \I__12293\ : InMux
    port map (
            O => \N__52690\,
            I => \N__52673\
        );

    \I__12292\ : InMux
    port map (
            O => \N__52689\,
            I => \N__52673\
        );

    \I__12291\ : InMux
    port map (
            O => \N__52688\,
            I => \N__52673\
        );

    \I__12290\ : InMux
    port map (
            O => \N__52687\,
            I => \N__52673\
        );

    \I__12289\ : LocalMux
    port map (
            O => \N__52684\,
            I => \N__52669\
        );

    \I__12288\ : LocalMux
    port map (
            O => \N__52673\,
            I => \N__52666\
        );

    \I__12287\ : InMux
    port map (
            O => \N__52672\,
            I => \N__52663\
        );

    \I__12286\ : Span4Mux_s1_h
    port map (
            O => \N__52669\,
            I => \N__52656\
        );

    \I__12285\ : Span4Mux_v
    port map (
            O => \N__52666\,
            I => \N__52656\
        );

    \I__12284\ : LocalMux
    port map (
            O => \N__52663\,
            I => \N__52656\
        );

    \I__12283\ : Span4Mux_h
    port map (
            O => \N__52656\,
            I => \N__52653\
        );

    \I__12282\ : Odrv4
    port map (
            O => \N__52653\,
            I => \current_shift_inst.PI_CTRL.N_150\
        );

    \I__12281\ : InMux
    port map (
            O => \N__52650\,
            I => \N__52635\
        );

    \I__12280\ : InMux
    port map (
            O => \N__52649\,
            I => \N__52635\
        );

    \I__12279\ : InMux
    port map (
            O => \N__52648\,
            I => \N__52635\
        );

    \I__12278\ : InMux
    port map (
            O => \N__52647\,
            I => \N__52635\
        );

    \I__12277\ : InMux
    port map (
            O => \N__52646\,
            I => \N__52635\
        );

    \I__12276\ : LocalMux
    port map (
            O => \N__52635\,
            I => \N__52631\
        );

    \I__12275\ : InMux
    port map (
            O => \N__52634\,
            I => \N__52628\
        );

    \I__12274\ : Span4Mux_v
    port map (
            O => \N__52631\,
            I => \N__52621\
        );

    \I__12273\ : LocalMux
    port map (
            O => \N__52628\,
            I => \N__52618\
        );

    \I__12272\ : InMux
    port map (
            O => \N__52627\,
            I => \N__52609\
        );

    \I__12271\ : InMux
    port map (
            O => \N__52626\,
            I => \N__52609\
        );

    \I__12270\ : InMux
    port map (
            O => \N__52625\,
            I => \N__52609\
        );

    \I__12269\ : InMux
    port map (
            O => \N__52624\,
            I => \N__52609\
        );

    \I__12268\ : Span4Mux_h
    port map (
            O => \N__52621\,
            I => \N__52606\
        );

    \I__12267\ : Span4Mux_v
    port map (
            O => \N__52618\,
            I => \N__52603\
        );

    \I__12266\ : LocalMux
    port map (
            O => \N__52609\,
            I => \N__52600\
        );

    \I__12265\ : Sp12to4
    port map (
            O => \N__52606\,
            I => \N__52593\
        );

    \I__12264\ : Sp12to4
    port map (
            O => \N__52603\,
            I => \N__52593\
        );

    \I__12263\ : Span12Mux_s4_h
    port map (
            O => \N__52600\,
            I => \N__52593\
        );

    \I__12262\ : Odrv12
    port map (
            O => \N__52593\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__12261\ : CascadeMux
    port map (
            O => \N__52590\,
            I => \N__52583\
        );

    \I__12260\ : CascadeMux
    port map (
            O => \N__52589\,
            I => \N__52580\
        );

    \I__12259\ : CascadeMux
    port map (
            O => \N__52588\,
            I => \N__52577\
        );

    \I__12258\ : InMux
    port map (
            O => \N__52587\,
            I => \N__52566\
        );

    \I__12257\ : InMux
    port map (
            O => \N__52586\,
            I => \N__52566\
        );

    \I__12256\ : InMux
    port map (
            O => \N__52583\,
            I => \N__52566\
        );

    \I__12255\ : InMux
    port map (
            O => \N__52580\,
            I => \N__52566\
        );

    \I__12254\ : InMux
    port map (
            O => \N__52577\,
            I => \N__52566\
        );

    \I__12253\ : LocalMux
    port map (
            O => \N__52566\,
            I => \N__52563\
        );

    \I__12252\ : Span4Mux_v
    port map (
            O => \N__52563\,
            I => \N__52557\
        );

    \I__12251\ : InMux
    port map (
            O => \N__52562\,
            I => \N__52552\
        );

    \I__12250\ : InMux
    port map (
            O => \N__52561\,
            I => \N__52552\
        );

    \I__12249\ : InMux
    port map (
            O => \N__52560\,
            I => \N__52549\
        );

    \I__12248\ : Sp12to4
    port map (
            O => \N__52557\,
            I => \N__52542\
        );

    \I__12247\ : LocalMux
    port map (
            O => \N__52552\,
            I => \N__52542\
        );

    \I__12246\ : LocalMux
    port map (
            O => \N__52549\,
            I => \N__52542\
        );

    \I__12245\ : Span12Mux_s9_h
    port map (
            O => \N__52542\,
            I => \N__52539\
        );

    \I__12244\ : Odrv12
    port map (
            O => \N__52539\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_11\
        );

    \I__12243\ : InMux
    port map (
            O => \N__52536\,
            I => \N__52533\
        );

    \I__12242\ : LocalMux
    port map (
            O => \N__52533\,
            I => \N__52528\
        );

    \I__12241\ : InMux
    port map (
            O => \N__52532\,
            I => \N__52523\
        );

    \I__12240\ : InMux
    port map (
            O => \N__52531\,
            I => \N__52523\
        );

    \I__12239\ : Span4Mux_s3_h
    port map (
            O => \N__52528\,
            I => \N__52518\
        );

    \I__12238\ : LocalMux
    port map (
            O => \N__52523\,
            I => \N__52518\
        );

    \I__12237\ : Span4Mux_v
    port map (
            O => \N__52518\,
            I => \N__52515\
        );

    \I__12236\ : Sp12to4
    port map (
            O => \N__52515\,
            I => \N__52512\
        );

    \I__12235\ : Odrv12
    port map (
            O => \N__52512\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__12234\ : InMux
    port map (
            O => \N__52509\,
            I => \N__52506\
        );

    \I__12233\ : LocalMux
    port map (
            O => \N__52506\,
            I => \N__52503\
        );

    \I__12232\ : Odrv4
    port map (
            O => \N__52503\,
            I => pwm_duty_input_7
        );

    \I__12231\ : ClkMux
    port map (
            O => \N__52500\,
            I => \N__52092\
        );

    \I__12230\ : ClkMux
    port map (
            O => \N__52499\,
            I => \N__52092\
        );

    \I__12229\ : ClkMux
    port map (
            O => \N__52498\,
            I => \N__52092\
        );

    \I__12228\ : ClkMux
    port map (
            O => \N__52497\,
            I => \N__52092\
        );

    \I__12227\ : ClkMux
    port map (
            O => \N__52496\,
            I => \N__52092\
        );

    \I__12226\ : ClkMux
    port map (
            O => \N__52495\,
            I => \N__52092\
        );

    \I__12225\ : ClkMux
    port map (
            O => \N__52494\,
            I => \N__52092\
        );

    \I__12224\ : ClkMux
    port map (
            O => \N__52493\,
            I => \N__52092\
        );

    \I__12223\ : ClkMux
    port map (
            O => \N__52492\,
            I => \N__52092\
        );

    \I__12222\ : ClkMux
    port map (
            O => \N__52491\,
            I => \N__52092\
        );

    \I__12221\ : ClkMux
    port map (
            O => \N__52490\,
            I => \N__52092\
        );

    \I__12220\ : ClkMux
    port map (
            O => \N__52489\,
            I => \N__52092\
        );

    \I__12219\ : ClkMux
    port map (
            O => \N__52488\,
            I => \N__52092\
        );

    \I__12218\ : ClkMux
    port map (
            O => \N__52487\,
            I => \N__52092\
        );

    \I__12217\ : ClkMux
    port map (
            O => \N__52486\,
            I => \N__52092\
        );

    \I__12216\ : ClkMux
    port map (
            O => \N__52485\,
            I => \N__52092\
        );

    \I__12215\ : ClkMux
    port map (
            O => \N__52484\,
            I => \N__52092\
        );

    \I__12214\ : ClkMux
    port map (
            O => \N__52483\,
            I => \N__52092\
        );

    \I__12213\ : ClkMux
    port map (
            O => \N__52482\,
            I => \N__52092\
        );

    \I__12212\ : ClkMux
    port map (
            O => \N__52481\,
            I => \N__52092\
        );

    \I__12211\ : ClkMux
    port map (
            O => \N__52480\,
            I => \N__52092\
        );

    \I__12210\ : ClkMux
    port map (
            O => \N__52479\,
            I => \N__52092\
        );

    \I__12209\ : ClkMux
    port map (
            O => \N__52478\,
            I => \N__52092\
        );

    \I__12208\ : ClkMux
    port map (
            O => \N__52477\,
            I => \N__52092\
        );

    \I__12207\ : ClkMux
    port map (
            O => \N__52476\,
            I => \N__52092\
        );

    \I__12206\ : ClkMux
    port map (
            O => \N__52475\,
            I => \N__52092\
        );

    \I__12205\ : ClkMux
    port map (
            O => \N__52474\,
            I => \N__52092\
        );

    \I__12204\ : ClkMux
    port map (
            O => \N__52473\,
            I => \N__52092\
        );

    \I__12203\ : ClkMux
    port map (
            O => \N__52472\,
            I => \N__52092\
        );

    \I__12202\ : ClkMux
    port map (
            O => \N__52471\,
            I => \N__52092\
        );

    \I__12201\ : ClkMux
    port map (
            O => \N__52470\,
            I => \N__52092\
        );

    \I__12200\ : ClkMux
    port map (
            O => \N__52469\,
            I => \N__52092\
        );

    \I__12199\ : ClkMux
    port map (
            O => \N__52468\,
            I => \N__52092\
        );

    \I__12198\ : ClkMux
    port map (
            O => \N__52467\,
            I => \N__52092\
        );

    \I__12197\ : ClkMux
    port map (
            O => \N__52466\,
            I => \N__52092\
        );

    \I__12196\ : ClkMux
    port map (
            O => \N__52465\,
            I => \N__52092\
        );

    \I__12195\ : ClkMux
    port map (
            O => \N__52464\,
            I => \N__52092\
        );

    \I__12194\ : ClkMux
    port map (
            O => \N__52463\,
            I => \N__52092\
        );

    \I__12193\ : ClkMux
    port map (
            O => \N__52462\,
            I => \N__52092\
        );

    \I__12192\ : ClkMux
    port map (
            O => \N__52461\,
            I => \N__52092\
        );

    \I__12191\ : ClkMux
    port map (
            O => \N__52460\,
            I => \N__52092\
        );

    \I__12190\ : ClkMux
    port map (
            O => \N__52459\,
            I => \N__52092\
        );

    \I__12189\ : ClkMux
    port map (
            O => \N__52458\,
            I => \N__52092\
        );

    \I__12188\ : ClkMux
    port map (
            O => \N__52457\,
            I => \N__52092\
        );

    \I__12187\ : ClkMux
    port map (
            O => \N__52456\,
            I => \N__52092\
        );

    \I__12186\ : ClkMux
    port map (
            O => \N__52455\,
            I => \N__52092\
        );

    \I__12185\ : ClkMux
    port map (
            O => \N__52454\,
            I => \N__52092\
        );

    \I__12184\ : ClkMux
    port map (
            O => \N__52453\,
            I => \N__52092\
        );

    \I__12183\ : ClkMux
    port map (
            O => \N__52452\,
            I => \N__52092\
        );

    \I__12182\ : ClkMux
    port map (
            O => \N__52451\,
            I => \N__52092\
        );

    \I__12181\ : ClkMux
    port map (
            O => \N__52450\,
            I => \N__52092\
        );

    \I__12180\ : ClkMux
    port map (
            O => \N__52449\,
            I => \N__52092\
        );

    \I__12179\ : ClkMux
    port map (
            O => \N__52448\,
            I => \N__52092\
        );

    \I__12178\ : ClkMux
    port map (
            O => \N__52447\,
            I => \N__52092\
        );

    \I__12177\ : ClkMux
    port map (
            O => \N__52446\,
            I => \N__52092\
        );

    \I__12176\ : ClkMux
    port map (
            O => \N__52445\,
            I => \N__52092\
        );

    \I__12175\ : ClkMux
    port map (
            O => \N__52444\,
            I => \N__52092\
        );

    \I__12174\ : ClkMux
    port map (
            O => \N__52443\,
            I => \N__52092\
        );

    \I__12173\ : ClkMux
    port map (
            O => \N__52442\,
            I => \N__52092\
        );

    \I__12172\ : ClkMux
    port map (
            O => \N__52441\,
            I => \N__52092\
        );

    \I__12171\ : ClkMux
    port map (
            O => \N__52440\,
            I => \N__52092\
        );

    \I__12170\ : ClkMux
    port map (
            O => \N__52439\,
            I => \N__52092\
        );

    \I__12169\ : ClkMux
    port map (
            O => \N__52438\,
            I => \N__52092\
        );

    \I__12168\ : ClkMux
    port map (
            O => \N__52437\,
            I => \N__52092\
        );

    \I__12167\ : ClkMux
    port map (
            O => \N__52436\,
            I => \N__52092\
        );

    \I__12166\ : ClkMux
    port map (
            O => \N__52435\,
            I => \N__52092\
        );

    \I__12165\ : ClkMux
    port map (
            O => \N__52434\,
            I => \N__52092\
        );

    \I__12164\ : ClkMux
    port map (
            O => \N__52433\,
            I => \N__52092\
        );

    \I__12163\ : ClkMux
    port map (
            O => \N__52432\,
            I => \N__52092\
        );

    \I__12162\ : ClkMux
    port map (
            O => \N__52431\,
            I => \N__52092\
        );

    \I__12161\ : ClkMux
    port map (
            O => \N__52430\,
            I => \N__52092\
        );

    \I__12160\ : ClkMux
    port map (
            O => \N__52429\,
            I => \N__52092\
        );

    \I__12159\ : ClkMux
    port map (
            O => \N__52428\,
            I => \N__52092\
        );

    \I__12158\ : ClkMux
    port map (
            O => \N__52427\,
            I => \N__52092\
        );

    \I__12157\ : ClkMux
    port map (
            O => \N__52426\,
            I => \N__52092\
        );

    \I__12156\ : ClkMux
    port map (
            O => \N__52425\,
            I => \N__52092\
        );

    \I__12155\ : ClkMux
    port map (
            O => \N__52424\,
            I => \N__52092\
        );

    \I__12154\ : ClkMux
    port map (
            O => \N__52423\,
            I => \N__52092\
        );

    \I__12153\ : ClkMux
    port map (
            O => \N__52422\,
            I => \N__52092\
        );

    \I__12152\ : ClkMux
    port map (
            O => \N__52421\,
            I => \N__52092\
        );

    \I__12151\ : ClkMux
    port map (
            O => \N__52420\,
            I => \N__52092\
        );

    \I__12150\ : ClkMux
    port map (
            O => \N__52419\,
            I => \N__52092\
        );

    \I__12149\ : ClkMux
    port map (
            O => \N__52418\,
            I => \N__52092\
        );

    \I__12148\ : ClkMux
    port map (
            O => \N__52417\,
            I => \N__52092\
        );

    \I__12147\ : ClkMux
    port map (
            O => \N__52416\,
            I => \N__52092\
        );

    \I__12146\ : ClkMux
    port map (
            O => \N__52415\,
            I => \N__52092\
        );

    \I__12145\ : ClkMux
    port map (
            O => \N__52414\,
            I => \N__52092\
        );

    \I__12144\ : ClkMux
    port map (
            O => \N__52413\,
            I => \N__52092\
        );

    \I__12143\ : ClkMux
    port map (
            O => \N__52412\,
            I => \N__52092\
        );

    \I__12142\ : ClkMux
    port map (
            O => \N__52411\,
            I => \N__52092\
        );

    \I__12141\ : ClkMux
    port map (
            O => \N__52410\,
            I => \N__52092\
        );

    \I__12140\ : ClkMux
    port map (
            O => \N__52409\,
            I => \N__52092\
        );

    \I__12139\ : ClkMux
    port map (
            O => \N__52408\,
            I => \N__52092\
        );

    \I__12138\ : ClkMux
    port map (
            O => \N__52407\,
            I => \N__52092\
        );

    \I__12137\ : ClkMux
    port map (
            O => \N__52406\,
            I => \N__52092\
        );

    \I__12136\ : ClkMux
    port map (
            O => \N__52405\,
            I => \N__52092\
        );

    \I__12135\ : ClkMux
    port map (
            O => \N__52404\,
            I => \N__52092\
        );

    \I__12134\ : ClkMux
    port map (
            O => \N__52403\,
            I => \N__52092\
        );

    \I__12133\ : ClkMux
    port map (
            O => \N__52402\,
            I => \N__52092\
        );

    \I__12132\ : ClkMux
    port map (
            O => \N__52401\,
            I => \N__52092\
        );

    \I__12131\ : ClkMux
    port map (
            O => \N__52400\,
            I => \N__52092\
        );

    \I__12130\ : ClkMux
    port map (
            O => \N__52399\,
            I => \N__52092\
        );

    \I__12129\ : ClkMux
    port map (
            O => \N__52398\,
            I => \N__52092\
        );

    \I__12128\ : ClkMux
    port map (
            O => \N__52397\,
            I => \N__52092\
        );

    \I__12127\ : ClkMux
    port map (
            O => \N__52396\,
            I => \N__52092\
        );

    \I__12126\ : ClkMux
    port map (
            O => \N__52395\,
            I => \N__52092\
        );

    \I__12125\ : ClkMux
    port map (
            O => \N__52394\,
            I => \N__52092\
        );

    \I__12124\ : ClkMux
    port map (
            O => \N__52393\,
            I => \N__52092\
        );

    \I__12123\ : ClkMux
    port map (
            O => \N__52392\,
            I => \N__52092\
        );

    \I__12122\ : ClkMux
    port map (
            O => \N__52391\,
            I => \N__52092\
        );

    \I__12121\ : ClkMux
    port map (
            O => \N__52390\,
            I => \N__52092\
        );

    \I__12120\ : ClkMux
    port map (
            O => \N__52389\,
            I => \N__52092\
        );

    \I__12119\ : ClkMux
    port map (
            O => \N__52388\,
            I => \N__52092\
        );

    \I__12118\ : ClkMux
    port map (
            O => \N__52387\,
            I => \N__52092\
        );

    \I__12117\ : ClkMux
    port map (
            O => \N__52386\,
            I => \N__52092\
        );

    \I__12116\ : ClkMux
    port map (
            O => \N__52385\,
            I => \N__52092\
        );

    \I__12115\ : ClkMux
    port map (
            O => \N__52384\,
            I => \N__52092\
        );

    \I__12114\ : ClkMux
    port map (
            O => \N__52383\,
            I => \N__52092\
        );

    \I__12113\ : ClkMux
    port map (
            O => \N__52382\,
            I => \N__52092\
        );

    \I__12112\ : ClkMux
    port map (
            O => \N__52381\,
            I => \N__52092\
        );

    \I__12111\ : ClkMux
    port map (
            O => \N__52380\,
            I => \N__52092\
        );

    \I__12110\ : ClkMux
    port map (
            O => \N__52379\,
            I => \N__52092\
        );

    \I__12109\ : ClkMux
    port map (
            O => \N__52378\,
            I => \N__52092\
        );

    \I__12108\ : ClkMux
    port map (
            O => \N__52377\,
            I => \N__52092\
        );

    \I__12107\ : ClkMux
    port map (
            O => \N__52376\,
            I => \N__52092\
        );

    \I__12106\ : ClkMux
    port map (
            O => \N__52375\,
            I => \N__52092\
        );

    \I__12105\ : ClkMux
    port map (
            O => \N__52374\,
            I => \N__52092\
        );

    \I__12104\ : ClkMux
    port map (
            O => \N__52373\,
            I => \N__52092\
        );

    \I__12103\ : ClkMux
    port map (
            O => \N__52372\,
            I => \N__52092\
        );

    \I__12102\ : ClkMux
    port map (
            O => \N__52371\,
            I => \N__52092\
        );

    \I__12101\ : ClkMux
    port map (
            O => \N__52370\,
            I => \N__52092\
        );

    \I__12100\ : ClkMux
    port map (
            O => \N__52369\,
            I => \N__52092\
        );

    \I__12099\ : ClkMux
    port map (
            O => \N__52368\,
            I => \N__52092\
        );

    \I__12098\ : ClkMux
    port map (
            O => \N__52367\,
            I => \N__52092\
        );

    \I__12097\ : ClkMux
    port map (
            O => \N__52366\,
            I => \N__52092\
        );

    \I__12096\ : ClkMux
    port map (
            O => \N__52365\,
            I => \N__52092\
        );

    \I__12095\ : GlobalMux
    port map (
            O => \N__52092\,
            I => clk_100mhz_0
        );

    \I__12094\ : InMux
    port map (
            O => \N__52089\,
            I => \N__52079\
        );

    \I__12093\ : InMux
    port map (
            O => \N__52088\,
            I => \N__52076\
        );

    \I__12092\ : InMux
    port map (
            O => \N__52087\,
            I => \N__52073\
        );

    \I__12091\ : InMux
    port map (
            O => \N__52086\,
            I => \N__52070\
        );

    \I__12090\ : InMux
    port map (
            O => \N__52085\,
            I => \N__52067\
        );

    \I__12089\ : InMux
    port map (
            O => \N__52084\,
            I => \N__52064\
        );

    \I__12088\ : InMux
    port map (
            O => \N__52083\,
            I => \N__52061\
        );

    \I__12087\ : InMux
    port map (
            O => \N__52082\,
            I => \N__52058\
        );

    \I__12086\ : LocalMux
    port map (
            O => \N__52079\,
            I => \N__52055\
        );

    \I__12085\ : LocalMux
    port map (
            O => \N__52076\,
            I => \N__52052\
        );

    \I__12084\ : LocalMux
    port map (
            O => \N__52073\,
            I => \N__52049\
        );

    \I__12083\ : LocalMux
    port map (
            O => \N__52070\,
            I => \N__52027\
        );

    \I__12082\ : LocalMux
    port map (
            O => \N__52067\,
            I => \N__51983\
        );

    \I__12081\ : LocalMux
    port map (
            O => \N__52064\,
            I => \N__51948\
        );

    \I__12080\ : LocalMux
    port map (
            O => \N__52061\,
            I => \N__51936\
        );

    \I__12079\ : LocalMux
    port map (
            O => \N__52058\,
            I => \N__51929\
        );

    \I__12078\ : Glb2LocalMux
    port map (
            O => \N__52055\,
            I => \N__51699\
        );

    \I__12077\ : Glb2LocalMux
    port map (
            O => \N__52052\,
            I => \N__51699\
        );

    \I__12076\ : Glb2LocalMux
    port map (
            O => \N__52049\,
            I => \N__51699\
        );

    \I__12075\ : SRMux
    port map (
            O => \N__52048\,
            I => \N__51699\
        );

    \I__12074\ : SRMux
    port map (
            O => \N__52047\,
            I => \N__51699\
        );

    \I__12073\ : SRMux
    port map (
            O => \N__52046\,
            I => \N__51699\
        );

    \I__12072\ : SRMux
    port map (
            O => \N__52045\,
            I => \N__51699\
        );

    \I__12071\ : SRMux
    port map (
            O => \N__52044\,
            I => \N__51699\
        );

    \I__12070\ : SRMux
    port map (
            O => \N__52043\,
            I => \N__51699\
        );

    \I__12069\ : SRMux
    port map (
            O => \N__52042\,
            I => \N__51699\
        );

    \I__12068\ : SRMux
    port map (
            O => \N__52041\,
            I => \N__51699\
        );

    \I__12067\ : SRMux
    port map (
            O => \N__52040\,
            I => \N__51699\
        );

    \I__12066\ : SRMux
    port map (
            O => \N__52039\,
            I => \N__51699\
        );

    \I__12065\ : SRMux
    port map (
            O => \N__52038\,
            I => \N__51699\
        );

    \I__12064\ : SRMux
    port map (
            O => \N__52037\,
            I => \N__51699\
        );

    \I__12063\ : SRMux
    port map (
            O => \N__52036\,
            I => \N__51699\
        );

    \I__12062\ : SRMux
    port map (
            O => \N__52035\,
            I => \N__51699\
        );

    \I__12061\ : SRMux
    port map (
            O => \N__52034\,
            I => \N__51699\
        );

    \I__12060\ : SRMux
    port map (
            O => \N__52033\,
            I => \N__51699\
        );

    \I__12059\ : SRMux
    port map (
            O => \N__52032\,
            I => \N__51699\
        );

    \I__12058\ : SRMux
    port map (
            O => \N__52031\,
            I => \N__51699\
        );

    \I__12057\ : SRMux
    port map (
            O => \N__52030\,
            I => \N__51699\
        );

    \I__12056\ : Glb2LocalMux
    port map (
            O => \N__52027\,
            I => \N__51699\
        );

    \I__12055\ : SRMux
    port map (
            O => \N__52026\,
            I => \N__51699\
        );

    \I__12054\ : SRMux
    port map (
            O => \N__52025\,
            I => \N__51699\
        );

    \I__12053\ : SRMux
    port map (
            O => \N__52024\,
            I => \N__51699\
        );

    \I__12052\ : SRMux
    port map (
            O => \N__52023\,
            I => \N__51699\
        );

    \I__12051\ : SRMux
    port map (
            O => \N__52022\,
            I => \N__51699\
        );

    \I__12050\ : SRMux
    port map (
            O => \N__52021\,
            I => \N__51699\
        );

    \I__12049\ : SRMux
    port map (
            O => \N__52020\,
            I => \N__51699\
        );

    \I__12048\ : SRMux
    port map (
            O => \N__52019\,
            I => \N__51699\
        );

    \I__12047\ : SRMux
    port map (
            O => \N__52018\,
            I => \N__51699\
        );

    \I__12046\ : SRMux
    port map (
            O => \N__52017\,
            I => \N__51699\
        );

    \I__12045\ : SRMux
    port map (
            O => \N__52016\,
            I => \N__51699\
        );

    \I__12044\ : SRMux
    port map (
            O => \N__52015\,
            I => \N__51699\
        );

    \I__12043\ : SRMux
    port map (
            O => \N__52014\,
            I => \N__51699\
        );

    \I__12042\ : SRMux
    port map (
            O => \N__52013\,
            I => \N__51699\
        );

    \I__12041\ : SRMux
    port map (
            O => \N__52012\,
            I => \N__51699\
        );

    \I__12040\ : SRMux
    port map (
            O => \N__52011\,
            I => \N__51699\
        );

    \I__12039\ : SRMux
    port map (
            O => \N__52010\,
            I => \N__51699\
        );

    \I__12038\ : SRMux
    port map (
            O => \N__52009\,
            I => \N__51699\
        );

    \I__12037\ : SRMux
    port map (
            O => \N__52008\,
            I => \N__51699\
        );

    \I__12036\ : SRMux
    port map (
            O => \N__52007\,
            I => \N__51699\
        );

    \I__12035\ : SRMux
    port map (
            O => \N__52006\,
            I => \N__51699\
        );

    \I__12034\ : SRMux
    port map (
            O => \N__52005\,
            I => \N__51699\
        );

    \I__12033\ : SRMux
    port map (
            O => \N__52004\,
            I => \N__51699\
        );

    \I__12032\ : SRMux
    port map (
            O => \N__52003\,
            I => \N__51699\
        );

    \I__12031\ : SRMux
    port map (
            O => \N__52002\,
            I => \N__51699\
        );

    \I__12030\ : SRMux
    port map (
            O => \N__52001\,
            I => \N__51699\
        );

    \I__12029\ : SRMux
    port map (
            O => \N__52000\,
            I => \N__51699\
        );

    \I__12028\ : SRMux
    port map (
            O => \N__51999\,
            I => \N__51699\
        );

    \I__12027\ : SRMux
    port map (
            O => \N__51998\,
            I => \N__51699\
        );

    \I__12026\ : SRMux
    port map (
            O => \N__51997\,
            I => \N__51699\
        );

    \I__12025\ : SRMux
    port map (
            O => \N__51996\,
            I => \N__51699\
        );

    \I__12024\ : SRMux
    port map (
            O => \N__51995\,
            I => \N__51699\
        );

    \I__12023\ : SRMux
    port map (
            O => \N__51994\,
            I => \N__51699\
        );

    \I__12022\ : SRMux
    port map (
            O => \N__51993\,
            I => \N__51699\
        );

    \I__12021\ : SRMux
    port map (
            O => \N__51992\,
            I => \N__51699\
        );

    \I__12020\ : SRMux
    port map (
            O => \N__51991\,
            I => \N__51699\
        );

    \I__12019\ : SRMux
    port map (
            O => \N__51990\,
            I => \N__51699\
        );

    \I__12018\ : SRMux
    port map (
            O => \N__51989\,
            I => \N__51699\
        );

    \I__12017\ : SRMux
    port map (
            O => \N__51988\,
            I => \N__51699\
        );

    \I__12016\ : SRMux
    port map (
            O => \N__51987\,
            I => \N__51699\
        );

    \I__12015\ : SRMux
    port map (
            O => \N__51986\,
            I => \N__51699\
        );

    \I__12014\ : Glb2LocalMux
    port map (
            O => \N__51983\,
            I => \N__51699\
        );

    \I__12013\ : SRMux
    port map (
            O => \N__51982\,
            I => \N__51699\
        );

    \I__12012\ : SRMux
    port map (
            O => \N__51981\,
            I => \N__51699\
        );

    \I__12011\ : SRMux
    port map (
            O => \N__51980\,
            I => \N__51699\
        );

    \I__12010\ : SRMux
    port map (
            O => \N__51979\,
            I => \N__51699\
        );

    \I__12009\ : SRMux
    port map (
            O => \N__51978\,
            I => \N__51699\
        );

    \I__12008\ : SRMux
    port map (
            O => \N__51977\,
            I => \N__51699\
        );

    \I__12007\ : SRMux
    port map (
            O => \N__51976\,
            I => \N__51699\
        );

    \I__12006\ : SRMux
    port map (
            O => \N__51975\,
            I => \N__51699\
        );

    \I__12005\ : SRMux
    port map (
            O => \N__51974\,
            I => \N__51699\
        );

    \I__12004\ : SRMux
    port map (
            O => \N__51973\,
            I => \N__51699\
        );

    \I__12003\ : SRMux
    port map (
            O => \N__51972\,
            I => \N__51699\
        );

    \I__12002\ : SRMux
    port map (
            O => \N__51971\,
            I => \N__51699\
        );

    \I__12001\ : SRMux
    port map (
            O => \N__51970\,
            I => \N__51699\
        );

    \I__12000\ : SRMux
    port map (
            O => \N__51969\,
            I => \N__51699\
        );

    \I__11999\ : SRMux
    port map (
            O => \N__51968\,
            I => \N__51699\
        );

    \I__11998\ : SRMux
    port map (
            O => \N__51967\,
            I => \N__51699\
        );

    \I__11997\ : SRMux
    port map (
            O => \N__51966\,
            I => \N__51699\
        );

    \I__11996\ : SRMux
    port map (
            O => \N__51965\,
            I => \N__51699\
        );

    \I__11995\ : SRMux
    port map (
            O => \N__51964\,
            I => \N__51699\
        );

    \I__11994\ : SRMux
    port map (
            O => \N__51963\,
            I => \N__51699\
        );

    \I__11993\ : SRMux
    port map (
            O => \N__51962\,
            I => \N__51699\
        );

    \I__11992\ : SRMux
    port map (
            O => \N__51961\,
            I => \N__51699\
        );

    \I__11991\ : SRMux
    port map (
            O => \N__51960\,
            I => \N__51699\
        );

    \I__11990\ : SRMux
    port map (
            O => \N__51959\,
            I => \N__51699\
        );

    \I__11989\ : SRMux
    port map (
            O => \N__51958\,
            I => \N__51699\
        );

    \I__11988\ : SRMux
    port map (
            O => \N__51957\,
            I => \N__51699\
        );

    \I__11987\ : SRMux
    port map (
            O => \N__51956\,
            I => \N__51699\
        );

    \I__11986\ : SRMux
    port map (
            O => \N__51955\,
            I => \N__51699\
        );

    \I__11985\ : SRMux
    port map (
            O => \N__51954\,
            I => \N__51699\
        );

    \I__11984\ : SRMux
    port map (
            O => \N__51953\,
            I => \N__51699\
        );

    \I__11983\ : SRMux
    port map (
            O => \N__51952\,
            I => \N__51699\
        );

    \I__11982\ : SRMux
    port map (
            O => \N__51951\,
            I => \N__51699\
        );

    \I__11981\ : Glb2LocalMux
    port map (
            O => \N__51948\,
            I => \N__51699\
        );

    \I__11980\ : SRMux
    port map (
            O => \N__51947\,
            I => \N__51699\
        );

    \I__11979\ : SRMux
    port map (
            O => \N__51946\,
            I => \N__51699\
        );

    \I__11978\ : SRMux
    port map (
            O => \N__51945\,
            I => \N__51699\
        );

    \I__11977\ : SRMux
    port map (
            O => \N__51944\,
            I => \N__51699\
        );

    \I__11976\ : SRMux
    port map (
            O => \N__51943\,
            I => \N__51699\
        );

    \I__11975\ : SRMux
    port map (
            O => \N__51942\,
            I => \N__51699\
        );

    \I__11974\ : SRMux
    port map (
            O => \N__51941\,
            I => \N__51699\
        );

    \I__11973\ : SRMux
    port map (
            O => \N__51940\,
            I => \N__51699\
        );

    \I__11972\ : SRMux
    port map (
            O => \N__51939\,
            I => \N__51699\
        );

    \I__11971\ : Glb2LocalMux
    port map (
            O => \N__51936\,
            I => \N__51699\
        );

    \I__11970\ : SRMux
    port map (
            O => \N__51935\,
            I => \N__51699\
        );

    \I__11969\ : SRMux
    port map (
            O => \N__51934\,
            I => \N__51699\
        );

    \I__11968\ : SRMux
    port map (
            O => \N__51933\,
            I => \N__51699\
        );

    \I__11967\ : SRMux
    port map (
            O => \N__51932\,
            I => \N__51699\
        );

    \I__11966\ : Glb2LocalMux
    port map (
            O => \N__51929\,
            I => \N__51699\
        );

    \I__11965\ : SRMux
    port map (
            O => \N__51928\,
            I => \N__51699\
        );

    \I__11964\ : GlobalMux
    port map (
            O => \N__51699\,
            I => \N__51696\
        );

    \I__11963\ : gio2CtrlBuf
    port map (
            O => \N__51696\,
            I => red_c_g
        );

    \I__11962\ : InMux
    port map (
            O => \N__51693\,
            I => \N__51690\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__51690\,
            I => \current_shift_inst.PI_CTRL.N_98\
        );

    \I__11960\ : CascadeMux
    port map (
            O => \N__51687\,
            I => \current_shift_inst.PI_CTRL.N_96_cascade_\
        );

    \I__11959\ : InMux
    port map (
            O => \N__51684\,
            I => \N__51681\
        );

    \I__11958\ : LocalMux
    port map (
            O => \N__51681\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__11957\ : InMux
    port map (
            O => \N__51678\,
            I => \N__51669\
        );

    \I__11956\ : InMux
    port map (
            O => \N__51677\,
            I => \N__51669\
        );

    \I__11955\ : InMux
    port map (
            O => \N__51676\,
            I => \N__51669\
        );

    \I__11954\ : LocalMux
    port map (
            O => \N__51669\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__11953\ : InMux
    port map (
            O => \N__51666\,
            I => \N__51663\
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__51663\,
            I => \N__51660\
        );

    \I__11951\ : Span12Mux_v
    port map (
            O => \N__51660\,
            I => \N__51657\
        );

    \I__11950\ : Span12Mux_h
    port map (
            O => \N__51657\,
            I => \N__51654\
        );

    \I__11949\ : Odrv12
    port map (
            O => \N__51654\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__11948\ : InMux
    port map (
            O => \N__51651\,
            I => \N__51648\
        );

    \I__11947\ : LocalMux
    port map (
            O => \N__51648\,
            I => \N__51645\
        );

    \I__11946\ : Span4Mux_v
    port map (
            O => \N__51645\,
            I => \N__51642\
        );

    \I__11945\ : Span4Mux_h
    port map (
            O => \N__51642\,
            I => \N__51639\
        );

    \I__11944\ : Sp12to4
    port map (
            O => \N__51639\,
            I => \N__51636\
        );

    \I__11943\ : Odrv12
    port map (
            O => \N__51636\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__11942\ : InMux
    port map (
            O => \N__51633\,
            I => \N__51630\
        );

    \I__11941\ : LocalMux
    port map (
            O => \N__51630\,
            I => \N__51627\
        );

    \I__11940\ : Span4Mux_v
    port map (
            O => \N__51627\,
            I => \N__51624\
        );

    \I__11939\ : Odrv4
    port map (
            O => \N__51624\,
            I => pwm_duty_input_2
        );

    \I__11938\ : InMux
    port map (
            O => \N__51621\,
            I => \N__51618\
        );

    \I__11937\ : LocalMux
    port map (
            O => \N__51618\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__11936\ : InMux
    port map (
            O => \N__51615\,
            I => \N__51612\
        );

    \I__11935\ : LocalMux
    port map (
            O => \N__51612\,
            I => \N__51609\
        );

    \I__11934\ : Odrv4
    port map (
            O => \N__51609\,
            I => pwm_duty_input_0
        );

    \I__11933\ : InMux
    port map (
            O => \N__51606\,
            I => \N__51597\
        );

    \I__11932\ : InMux
    port map (
            O => \N__51605\,
            I => \N__51597\
        );

    \I__11931\ : InMux
    port map (
            O => \N__51604\,
            I => \N__51597\
        );

    \I__11930\ : LocalMux
    port map (
            O => \N__51597\,
            I => \current_shift_inst.PI_CTRL.N_152\
        );

    \I__11929\ : InMux
    port map (
            O => \N__51594\,
            I => \N__51591\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__51591\,
            I => \N__51588\
        );

    \I__11927\ : Span4Mux_v
    port map (
            O => \N__51588\,
            I => \N__51585\
        );

    \I__11926\ : Sp12to4
    port map (
            O => \N__51585\,
            I => \N__51582\
        );

    \I__11925\ : Span12Mux_h
    port map (
            O => \N__51582\,
            I => \N__51579\
        );

    \I__11924\ : Odrv12
    port map (
            O => \N__51579\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__11923\ : InMux
    port map (
            O => \N__51576\,
            I => \N__51573\
        );

    \I__11922\ : LocalMux
    port map (
            O => \N__51573\,
            I => \N__51570\
        );

    \I__11921\ : Odrv4
    port map (
            O => \N__51570\,
            I => pwm_duty_input_1
        );

    \I__11920\ : InMux
    port map (
            O => \N__51567\,
            I => \N__51564\
        );

    \I__11919\ : LocalMux
    port map (
            O => \N__51564\,
            I => \N__51559\
        );

    \I__11918\ : InMux
    port map (
            O => \N__51563\,
            I => \N__51556\
        );

    \I__11917\ : InMux
    port map (
            O => \N__51562\,
            I => \N__51553\
        );

    \I__11916\ : Span4Mux_v
    port map (
            O => \N__51559\,
            I => \N__51550\
        );

    \I__11915\ : LocalMux
    port map (
            O => \N__51556\,
            I => \N__51545\
        );

    \I__11914\ : LocalMux
    port map (
            O => \N__51553\,
            I => \N__51545\
        );

    \I__11913\ : Sp12to4
    port map (
            O => \N__51550\,
            I => \N__51542\
        );

    \I__11912\ : Span12Mux_v
    port map (
            O => \N__51545\,
            I => \N__51539\
        );

    \I__11911\ : Span12Mux_s8_h
    port map (
            O => \N__51542\,
            I => \N__51536\
        );

    \I__11910\ : Span12Mux_h
    port map (
            O => \N__51539\,
            I => \N__51533\
        );

    \I__11909\ : Odrv12
    port map (
            O => \N__51536\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__11908\ : Odrv12
    port map (
            O => \N__51533\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__11907\ : InMux
    port map (
            O => \N__51528\,
            I => \N__51524\
        );

    \I__11906\ : InMux
    port map (
            O => \N__51527\,
            I => \N__51521\
        );

    \I__11905\ : LocalMux
    port map (
            O => \N__51524\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__11904\ : LocalMux
    port map (
            O => \N__51521\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__11903\ : InMux
    port map (
            O => \N__51516\,
            I => \N__51513\
        );

    \I__11902\ : LocalMux
    port map (
            O => \N__51513\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__11901\ : InMux
    port map (
            O => \N__51510\,
            I => \N__51507\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__51507\,
            I => \N__51504\
        );

    \I__11899\ : Span4Mux_s0_h
    port map (
            O => \N__51504\,
            I => \N__51501\
        );

    \I__11898\ : Odrv4
    port map (
            O => \N__51501\,
            I => pwm_duty_input_3
        );

    \I__11897\ : CascadeMux
    port map (
            O => \N__51498\,
            I => \N__51493\
        );

    \I__11896\ : InMux
    port map (
            O => \N__51497\,
            I => \N__51490\
        );

    \I__11895\ : InMux
    port map (
            O => \N__51496\,
            I => \N__51487\
        );

    \I__11894\ : InMux
    port map (
            O => \N__51493\,
            I => \N__51484\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__51490\,
            I => \N__51481\
        );

    \I__11892\ : LocalMux
    port map (
            O => \N__51487\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__51484\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__11890\ : Odrv12
    port map (
            O => \N__51481\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__11889\ : InMux
    port map (
            O => \N__51474\,
            I => \N__51471\
        );

    \I__11888\ : LocalMux
    port map (
            O => \N__51471\,
            I => \N__51468\
        );

    \I__11887\ : Odrv4
    port map (
            O => \N__51468\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\
        );

    \I__11886\ : InMux
    port map (
            O => \N__51465\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17\
        );

    \I__11885\ : InMux
    port map (
            O => \N__51462\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18\
        );

    \I__11884\ : InMux
    port map (
            O => \N__51459\,
            I => \N__51456\
        );

    \I__11883\ : LocalMux
    port map (
            O => \N__51456\,
            I => \N__51453\
        );

    \I__11882\ : Odrv4
    port map (
            O => \N__51453\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\
        );

    \I__11881\ : InMux
    port map (
            O => \N__51450\,
            I => \N__51446\
        );

    \I__11880\ : InMux
    port map (
            O => \N__51449\,
            I => \N__51443\
        );

    \I__11879\ : LocalMux
    port map (
            O => \N__51446\,
            I => \N__51440\
        );

    \I__11878\ : LocalMux
    port map (
            O => \N__51443\,
            I => \N__51437\
        );

    \I__11877\ : Span12Mux_h
    port map (
            O => \N__51440\,
            I => \N__51434\
        );

    \I__11876\ : Span4Mux_v
    port map (
            O => \N__51437\,
            I => \N__51431\
        );

    \I__11875\ : Odrv12
    port map (
            O => \N__51434\,
            I => \pwm_generator_inst.O_10\
        );

    \I__11874\ : Odrv4
    port map (
            O => \N__51431\,
            I => \pwm_generator_inst.O_10\
        );

    \I__11873\ : InMux
    port map (
            O => \N__51426\,
            I => \N__51422\
        );

    \I__11872\ : InMux
    port map (
            O => \N__51425\,
            I => \N__51418\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__51422\,
            I => \N__51415\
        );

    \I__11870\ : InMux
    port map (
            O => \N__51421\,
            I => \N__51412\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__51418\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__11868\ : Odrv12
    port map (
            O => \N__51415\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__51412\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__11866\ : InMux
    port map (
            O => \N__51405\,
            I => \N__51402\
        );

    \I__11865\ : LocalMux
    port map (
            O => \N__51402\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4\
        );

    \I__11864\ : InMux
    port map (
            O => \N__51399\,
            I => \N__51396\
        );

    \I__11863\ : LocalMux
    port map (
            O => \N__51396\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\
        );

    \I__11862\ : InMux
    port map (
            O => \N__51393\,
            I => \N__51390\
        );

    \I__11861\ : LocalMux
    port map (
            O => \N__51390\,
            I => \N__51387\
        );

    \I__11860\ : Odrv12
    port map (
            O => \N__51387\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\
        );

    \I__11859\ : InMux
    port map (
            O => \N__51384\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9\
        );

    \I__11858\ : CascadeMux
    port map (
            O => \N__51381\,
            I => \N__51375\
        );

    \I__11857\ : InMux
    port map (
            O => \N__51380\,
            I => \N__51371\
        );

    \I__11856\ : CascadeMux
    port map (
            O => \N__51379\,
            I => \N__51364\
        );

    \I__11855\ : CascadeMux
    port map (
            O => \N__51378\,
            I => \N__51361\
        );

    \I__11854\ : InMux
    port map (
            O => \N__51375\,
            I => \N__51355\
        );

    \I__11853\ : InMux
    port map (
            O => \N__51374\,
            I => \N__51352\
        );

    \I__11852\ : LocalMux
    port map (
            O => \N__51371\,
            I => \N__51349\
        );

    \I__11851\ : InMux
    port map (
            O => \N__51370\,
            I => \N__51346\
        );

    \I__11850\ : InMux
    port map (
            O => \N__51369\,
            I => \N__51337\
        );

    \I__11849\ : InMux
    port map (
            O => \N__51368\,
            I => \N__51337\
        );

    \I__11848\ : InMux
    port map (
            O => \N__51367\,
            I => \N__51337\
        );

    \I__11847\ : InMux
    port map (
            O => \N__51364\,
            I => \N__51337\
        );

    \I__11846\ : InMux
    port map (
            O => \N__51361\,
            I => \N__51328\
        );

    \I__11845\ : InMux
    port map (
            O => \N__51360\,
            I => \N__51328\
        );

    \I__11844\ : InMux
    port map (
            O => \N__51359\,
            I => \N__51328\
        );

    \I__11843\ : InMux
    port map (
            O => \N__51358\,
            I => \N__51328\
        );

    \I__11842\ : LocalMux
    port map (
            O => \N__51355\,
            I => \N__51323\
        );

    \I__11841\ : LocalMux
    port map (
            O => \N__51352\,
            I => \N__51323\
        );

    \I__11840\ : Span4Mux_h
    port map (
            O => \N__51349\,
            I => \N__51320\
        );

    \I__11839\ : LocalMux
    port map (
            O => \N__51346\,
            I => \N__51317\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__51337\,
            I => \N__51314\
        );

    \I__11837\ : LocalMux
    port map (
            O => \N__51328\,
            I => \N__51309\
        );

    \I__11836\ : Span4Mux_h
    port map (
            O => \N__51323\,
            I => \N__51309\
        );

    \I__11835\ : Odrv4
    port map (
            O => \N__51320\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__11834\ : Odrv12
    port map (
            O => \N__51317\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__11833\ : Odrv12
    port map (
            O => \N__51314\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__11832\ : Odrv4
    port map (
            O => \N__51309\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__11831\ : InMux
    port map (
            O => \N__51300\,
            I => \N__51296\
        );

    \I__11830\ : InMux
    port map (
            O => \N__51299\,
            I => \N__51293\
        );

    \I__11829\ : LocalMux
    port map (
            O => \N__51296\,
            I => \N__51290\
        );

    \I__11828\ : LocalMux
    port map (
            O => \N__51293\,
            I => \N__51287\
        );

    \I__11827\ : Span4Mux_v
    port map (
            O => \N__51290\,
            I => \N__51284\
        );

    \I__11826\ : Span4Mux_v
    port map (
            O => \N__51287\,
            I => \N__51279\
        );

    \I__11825\ : Span4Mux_h
    port map (
            O => \N__51284\,
            I => \N__51279\
        );

    \I__11824\ : Span4Mux_h
    port map (
            O => \N__51279\,
            I => \N__51276\
        );

    \I__11823\ : Odrv4
    port map (
            O => \N__51276\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__11822\ : InMux
    port map (
            O => \N__51273\,
            I => \N__51270\
        );

    \I__11821\ : LocalMux
    port map (
            O => \N__51270\,
            I => \N__51267\
        );

    \I__11820\ : Odrv4
    port map (
            O => \N__51267\,
            I => \pwm_generator_inst.un19_threshold_0_axb_1\
        );

    \I__11819\ : InMux
    port map (
            O => \N__51264\,
            I => \pwm_generator_inst.un15_threshold_1_cry_10\
        );

    \I__11818\ : InMux
    port map (
            O => \N__51261\,
            I => \N__51257\
        );

    \I__11817\ : InMux
    port map (
            O => \N__51260\,
            I => \N__51254\
        );

    \I__11816\ : LocalMux
    port map (
            O => \N__51257\,
            I => \N__51250\
        );

    \I__11815\ : LocalMux
    port map (
            O => \N__51254\,
            I => \N__51247\
        );

    \I__11814\ : InMux
    port map (
            O => \N__51253\,
            I => \N__51244\
        );

    \I__11813\ : Span4Mux_v
    port map (
            O => \N__51250\,
            I => \N__51239\
        );

    \I__11812\ : Span4Mux_h
    port map (
            O => \N__51247\,
            I => \N__51239\
        );

    \I__11811\ : LocalMux
    port map (
            O => \N__51244\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__11810\ : Odrv4
    port map (
            O => \N__51239\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__11809\ : InMux
    port map (
            O => \N__51234\,
            I => \N__51231\
        );

    \I__11808\ : LocalMux
    port map (
            O => \N__51231\,
            I => \N__51228\
        );

    \I__11807\ : Odrv12
    port map (
            O => \N__51228\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\
        );

    \I__11806\ : InMux
    port map (
            O => \N__51225\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11\
        );

    \I__11805\ : InMux
    port map (
            O => \N__51222\,
            I => \N__51218\
        );

    \I__11804\ : InMux
    port map (
            O => \N__51221\,
            I => \N__51215\
        );

    \I__11803\ : LocalMux
    port map (
            O => \N__51218\,
            I => \N__51212\
        );

    \I__11802\ : LocalMux
    port map (
            O => \N__51215\,
            I => \N__51207\
        );

    \I__11801\ : Span4Mux_h
    port map (
            O => \N__51212\,
            I => \N__51207\
        );

    \I__11800\ : Odrv4
    port map (
            O => \N__51207\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__11799\ : InMux
    port map (
            O => \N__51204\,
            I => \N__51201\
        );

    \I__11798\ : LocalMux
    port map (
            O => \N__51201\,
            I => \N__51198\
        );

    \I__11797\ : Odrv12
    port map (
            O => \N__51198\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\
        );

    \I__11796\ : InMux
    port map (
            O => \N__51195\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12\
        );

    \I__11795\ : InMux
    port map (
            O => \N__51192\,
            I => \N__51187\
        );

    \I__11794\ : InMux
    port map (
            O => \N__51191\,
            I => \N__51184\
        );

    \I__11793\ : InMux
    port map (
            O => \N__51190\,
            I => \N__51181\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__51187\,
            I => \N__51178\
        );

    \I__11791\ : LocalMux
    port map (
            O => \N__51184\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__11790\ : LocalMux
    port map (
            O => \N__51181\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__11789\ : Odrv12
    port map (
            O => \N__51178\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__11788\ : InMux
    port map (
            O => \N__51171\,
            I => \N__51168\
        );

    \I__11787\ : LocalMux
    port map (
            O => \N__51168\,
            I => \N__51165\
        );

    \I__11786\ : Span4Mux_h
    port map (
            O => \N__51165\,
            I => \N__51162\
        );

    \I__11785\ : Odrv4
    port map (
            O => \N__51162\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\
        );

    \I__11784\ : InMux
    port map (
            O => \N__51159\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13\
        );

    \I__11783\ : InMux
    port map (
            O => \N__51156\,
            I => \N__51153\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__51153\,
            I => \N__51150\
        );

    \I__11781\ : Span4Mux_h
    port map (
            O => \N__51150\,
            I => \N__51145\
        );

    \I__11780\ : InMux
    port map (
            O => \N__51149\,
            I => \N__51142\
        );

    \I__11779\ : InMux
    port map (
            O => \N__51148\,
            I => \N__51139\
        );

    \I__11778\ : Span4Mux_h
    port map (
            O => \N__51145\,
            I => \N__51136\
        );

    \I__11777\ : LocalMux
    port map (
            O => \N__51142\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__11776\ : LocalMux
    port map (
            O => \N__51139\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__11775\ : Odrv4
    port map (
            O => \N__51136\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__11774\ : InMux
    port map (
            O => \N__51129\,
            I => \N__51126\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__51126\,
            I => \N__51123\
        );

    \I__11772\ : Odrv12
    port map (
            O => \N__51123\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\
        );

    \I__11771\ : InMux
    port map (
            O => \N__51120\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14\
        );

    \I__11770\ : CascadeMux
    port map (
            O => \N__51117\,
            I => \N__51112\
        );

    \I__11769\ : InMux
    port map (
            O => \N__51116\,
            I => \N__51109\
        );

    \I__11768\ : InMux
    port map (
            O => \N__51115\,
            I => \N__51106\
        );

    \I__11767\ : InMux
    port map (
            O => \N__51112\,
            I => \N__51103\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__51109\,
            I => \N__51100\
        );

    \I__11765\ : LocalMux
    port map (
            O => \N__51106\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__51103\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__11763\ : Odrv12
    port map (
            O => \N__51100\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__11762\ : InMux
    port map (
            O => \N__51093\,
            I => \N__51090\
        );

    \I__11761\ : LocalMux
    port map (
            O => \N__51090\,
            I => \N__51087\
        );

    \I__11760\ : Odrv12
    port map (
            O => \N__51087\,
            I => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\
        );

    \I__11759\ : InMux
    port map (
            O => \N__51084\,
            I => \bfn_20_27_0_\
        );

    \I__11758\ : InMux
    port map (
            O => \N__51081\,
            I => \N__51077\
        );

    \I__11757\ : InMux
    port map (
            O => \N__51080\,
            I => \N__51074\
        );

    \I__11756\ : LocalMux
    port map (
            O => \N__51077\,
            I => \N__51071\
        );

    \I__11755\ : LocalMux
    port map (
            O => \N__51074\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__11754\ : Odrv12
    port map (
            O => \N__51071\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__11753\ : InMux
    port map (
            O => \N__51066\,
            I => \N__51063\
        );

    \I__11752\ : LocalMux
    port map (
            O => \N__51063\,
            I => \N__51060\
        );

    \I__11751\ : Span4Mux_h
    port map (
            O => \N__51060\,
            I => \N__51057\
        );

    \I__11750\ : Odrv4
    port map (
            O => \N__51057\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\
        );

    \I__11749\ : InMux
    port map (
            O => \N__51054\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16\
        );

    \I__11748\ : InMux
    port map (
            O => \N__51051\,
            I => \N__51048\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__51048\,
            I => \N__51045\
        );

    \I__11746\ : Span4Mux_v
    port map (
            O => \N__51045\,
            I => \N__51042\
        );

    \I__11745\ : Span4Mux_h
    port map (
            O => \N__51042\,
            I => \N__51039\
        );

    \I__11744\ : Odrv4
    port map (
            O => \N__51039\,
            I => \pwm_generator_inst.O_3\
        );

    \I__11743\ : InMux
    port map (
            O => \N__51036\,
            I => \N__51033\
        );

    \I__11742\ : LocalMux
    port map (
            O => \N__51033\,
            I => \pwm_generator_inst.un15_threshold_1_axb_3\
        );

    \I__11741\ : InMux
    port map (
            O => \N__51030\,
            I => \N__51027\
        );

    \I__11740\ : LocalMux
    port map (
            O => \N__51027\,
            I => \N__51024\
        );

    \I__11739\ : Span4Mux_v
    port map (
            O => \N__51024\,
            I => \N__51021\
        );

    \I__11738\ : Span4Mux_h
    port map (
            O => \N__51021\,
            I => \N__51018\
        );

    \I__11737\ : Odrv4
    port map (
            O => \N__51018\,
            I => \pwm_generator_inst.O_4\
        );

    \I__11736\ : InMux
    port map (
            O => \N__51015\,
            I => \N__51012\
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__51012\,
            I => \pwm_generator_inst.un15_threshold_1_axb_4\
        );

    \I__11734\ : InMux
    port map (
            O => \N__51009\,
            I => \N__51006\
        );

    \I__11733\ : LocalMux
    port map (
            O => \N__51006\,
            I => \N__51003\
        );

    \I__11732\ : Span4Mux_h
    port map (
            O => \N__51003\,
            I => \N__51000\
        );

    \I__11731\ : Span4Mux_h
    port map (
            O => \N__51000\,
            I => \N__50997\
        );

    \I__11730\ : Odrv4
    port map (
            O => \N__50997\,
            I => \pwm_generator_inst.O_5\
        );

    \I__11729\ : InMux
    port map (
            O => \N__50994\,
            I => \N__50991\
        );

    \I__11728\ : LocalMux
    port map (
            O => \N__50991\,
            I => \pwm_generator_inst.un15_threshold_1_axb_5\
        );

    \I__11727\ : InMux
    port map (
            O => \N__50988\,
            I => \N__50985\
        );

    \I__11726\ : LocalMux
    port map (
            O => \N__50985\,
            I => \N__50982\
        );

    \I__11725\ : Span4Mux_h
    port map (
            O => \N__50982\,
            I => \N__50979\
        );

    \I__11724\ : Span4Mux_h
    port map (
            O => \N__50979\,
            I => \N__50976\
        );

    \I__11723\ : Odrv4
    port map (
            O => \N__50976\,
            I => \pwm_generator_inst.O_6\
        );

    \I__11722\ : InMux
    port map (
            O => \N__50973\,
            I => \N__50970\
        );

    \I__11721\ : LocalMux
    port map (
            O => \N__50970\,
            I => \pwm_generator_inst.un15_threshold_1_axb_6\
        );

    \I__11720\ : InMux
    port map (
            O => \N__50967\,
            I => \N__50964\
        );

    \I__11719\ : LocalMux
    port map (
            O => \N__50964\,
            I => \N__50961\
        );

    \I__11718\ : Span4Mux_v
    port map (
            O => \N__50961\,
            I => \N__50958\
        );

    \I__11717\ : Span4Mux_h
    port map (
            O => \N__50958\,
            I => \N__50955\
        );

    \I__11716\ : Odrv4
    port map (
            O => \N__50955\,
            I => \pwm_generator_inst.O_7\
        );

    \I__11715\ : InMux
    port map (
            O => \N__50952\,
            I => \N__50949\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__50949\,
            I => \pwm_generator_inst.un15_threshold_1_axb_7\
        );

    \I__11713\ : InMux
    port map (
            O => \N__50946\,
            I => \N__50943\
        );

    \I__11712\ : LocalMux
    port map (
            O => \N__50943\,
            I => \N__50940\
        );

    \I__11711\ : Span4Mux_h
    port map (
            O => \N__50940\,
            I => \N__50937\
        );

    \I__11710\ : Span4Mux_h
    port map (
            O => \N__50937\,
            I => \N__50934\
        );

    \I__11709\ : Odrv4
    port map (
            O => \N__50934\,
            I => \pwm_generator_inst.O_8\
        );

    \I__11708\ : InMux
    port map (
            O => \N__50931\,
            I => \N__50928\
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__50928\,
            I => \pwm_generator_inst.un15_threshold_1_axb_8\
        );

    \I__11706\ : InMux
    port map (
            O => \N__50925\,
            I => \N__50922\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__50922\,
            I => \N__50919\
        );

    \I__11704\ : Span12Mux_s6_v
    port map (
            O => \N__50919\,
            I => \N__50916\
        );

    \I__11703\ : Odrv12
    port map (
            O => \N__50916\,
            I => \pwm_generator_inst.O_9\
        );

    \I__11702\ : InMux
    port map (
            O => \N__50913\,
            I => \N__50910\
        );

    \I__11701\ : LocalMux
    port map (
            O => \N__50910\,
            I => \pwm_generator_inst.un15_threshold_1_axb_9\
        );

    \I__11700\ : InMux
    port map (
            O => \N__50907\,
            I => \N__50904\
        );

    \I__11699\ : LocalMux
    port map (
            O => \N__50904\,
            I => \N__50901\
        );

    \I__11698\ : Odrv4
    port map (
            O => \N__50901\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\
        );

    \I__11697\ : InMux
    port map (
            O => \N__50898\,
            I => \N__50895\
        );

    \I__11696\ : LocalMux
    port map (
            O => \N__50895\,
            I => \N__50892\
        );

    \I__11695\ : Span4Mux_h
    port map (
            O => \N__50892\,
            I => \N__50888\
        );

    \I__11694\ : InMux
    port map (
            O => \N__50891\,
            I => \N__50885\
        );

    \I__11693\ : Odrv4
    port map (
            O => \N__50888\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__11692\ : LocalMux
    port map (
            O => \N__50885\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__11691\ : CascadeMux
    port map (
            O => \N__50880\,
            I => \N__50870\
        );

    \I__11690\ : InMux
    port map (
            O => \N__50879\,
            I => \N__50866\
        );

    \I__11689\ : InMux
    port map (
            O => \N__50878\,
            I => \N__50861\
        );

    \I__11688\ : InMux
    port map (
            O => \N__50877\,
            I => \N__50861\
        );

    \I__11687\ : InMux
    port map (
            O => \N__50876\,
            I => \N__50856\
        );

    \I__11686\ : InMux
    port map (
            O => \N__50875\,
            I => \N__50856\
        );

    \I__11685\ : InMux
    port map (
            O => \N__50874\,
            I => \N__50853\
        );

    \I__11684\ : InMux
    port map (
            O => \N__50873\,
            I => \N__50838\
        );

    \I__11683\ : InMux
    port map (
            O => \N__50870\,
            I => \N__50838\
        );

    \I__11682\ : InMux
    port map (
            O => \N__50869\,
            I => \N__50838\
        );

    \I__11681\ : LocalMux
    port map (
            O => \N__50866\,
            I => \N__50826\
        );

    \I__11680\ : LocalMux
    port map (
            O => \N__50861\,
            I => \N__50826\
        );

    \I__11679\ : LocalMux
    port map (
            O => \N__50856\,
            I => \N__50826\
        );

    \I__11678\ : LocalMux
    port map (
            O => \N__50853\,
            I => \N__50819\
        );

    \I__11677\ : InMux
    port map (
            O => \N__50852\,
            I => \N__50804\
        );

    \I__11676\ : InMux
    port map (
            O => \N__50851\,
            I => \N__50804\
        );

    \I__11675\ : InMux
    port map (
            O => \N__50850\,
            I => \N__50804\
        );

    \I__11674\ : InMux
    port map (
            O => \N__50849\,
            I => \N__50804\
        );

    \I__11673\ : InMux
    port map (
            O => \N__50848\,
            I => \N__50804\
        );

    \I__11672\ : InMux
    port map (
            O => \N__50847\,
            I => \N__50799\
        );

    \I__11671\ : InMux
    port map (
            O => \N__50846\,
            I => \N__50799\
        );

    \I__11670\ : InMux
    port map (
            O => \N__50845\,
            I => \N__50796\
        );

    \I__11669\ : LocalMux
    port map (
            O => \N__50838\,
            I => \N__50793\
        );

    \I__11668\ : InMux
    port map (
            O => \N__50837\,
            I => \N__50788\
        );

    \I__11667\ : InMux
    port map (
            O => \N__50836\,
            I => \N__50788\
        );

    \I__11666\ : InMux
    port map (
            O => \N__50835\,
            I => \N__50785\
        );

    \I__11665\ : InMux
    port map (
            O => \N__50834\,
            I => \N__50780\
        );

    \I__11664\ : InMux
    port map (
            O => \N__50833\,
            I => \N__50780\
        );

    \I__11663\ : Span4Mux_v
    port map (
            O => \N__50826\,
            I => \N__50777\
        );

    \I__11662\ : InMux
    port map (
            O => \N__50825\,
            I => \N__50768\
        );

    \I__11661\ : InMux
    port map (
            O => \N__50824\,
            I => \N__50768\
        );

    \I__11660\ : InMux
    port map (
            O => \N__50823\,
            I => \N__50768\
        );

    \I__11659\ : InMux
    port map (
            O => \N__50822\,
            I => \N__50768\
        );

    \I__11658\ : Span4Mux_h
    port map (
            O => \N__50819\,
            I => \N__50765\
        );

    \I__11657\ : InMux
    port map (
            O => \N__50818\,
            I => \N__50756\
        );

    \I__11656\ : InMux
    port map (
            O => \N__50817\,
            I => \N__50756\
        );

    \I__11655\ : InMux
    port map (
            O => \N__50816\,
            I => \N__50756\
        );

    \I__11654\ : InMux
    port map (
            O => \N__50815\,
            I => \N__50756\
        );

    \I__11653\ : LocalMux
    port map (
            O => \N__50804\,
            I => \N__50751\
        );

    \I__11652\ : LocalMux
    port map (
            O => \N__50799\,
            I => \N__50751\
        );

    \I__11651\ : LocalMux
    port map (
            O => \N__50796\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11650\ : Odrv4
    port map (
            O => \N__50793\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11649\ : LocalMux
    port map (
            O => \N__50788\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11648\ : LocalMux
    port map (
            O => \N__50785\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11647\ : LocalMux
    port map (
            O => \N__50780\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11646\ : Odrv4
    port map (
            O => \N__50777\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11645\ : LocalMux
    port map (
            O => \N__50768\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11644\ : Odrv4
    port map (
            O => \N__50765\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11643\ : LocalMux
    port map (
            O => \N__50756\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11642\ : Odrv4
    port map (
            O => \N__50751\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11641\ : InMux
    port map (
            O => \N__50730\,
            I => \N__50727\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__50727\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__11639\ : CascadeMux
    port map (
            O => \N__50724\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\
        );

    \I__11638\ : InMux
    port map (
            O => \N__50721\,
            I => \N__50718\
        );

    \I__11637\ : LocalMux
    port map (
            O => \N__50718\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29\
        );

    \I__11636\ : InMux
    port map (
            O => \N__50715\,
            I => \N__50712\
        );

    \I__11635\ : LocalMux
    port map (
            O => \N__50712\,
            I => \N__50709\
        );

    \I__11634\ : Span4Mux_h
    port map (
            O => \N__50709\,
            I => \N__50705\
        );

    \I__11633\ : InMux
    port map (
            O => \N__50708\,
            I => \N__50702\
        );

    \I__11632\ : Odrv4
    port map (
            O => \N__50705\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__11631\ : LocalMux
    port map (
            O => \N__50702\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__11630\ : InMux
    port map (
            O => \N__50697\,
            I => \N__50693\
        );

    \I__11629\ : CascadeMux
    port map (
            O => \N__50696\,
            I => \N__50690\
        );

    \I__11628\ : LocalMux
    port map (
            O => \N__50693\,
            I => \N__50687\
        );

    \I__11627\ : InMux
    port map (
            O => \N__50690\,
            I => \N__50684\
        );

    \I__11626\ : Odrv4
    port map (
            O => \N__50687\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__50684\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__11624\ : InMux
    port map (
            O => \N__50679\,
            I => \N__50676\
        );

    \I__11623\ : LocalMux
    port map (
            O => \N__50676\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\
        );

    \I__11622\ : CascadeMux
    port map (
            O => \N__50673\,
            I => \N__50669\
        );

    \I__11621\ : InMux
    port map (
            O => \N__50672\,
            I => \N__50666\
        );

    \I__11620\ : InMux
    port map (
            O => \N__50669\,
            I => \N__50663\
        );

    \I__11619\ : LocalMux
    port map (
            O => \N__50666\,
            I => \N__50657\
        );

    \I__11618\ : LocalMux
    port map (
            O => \N__50663\,
            I => \N__50657\
        );

    \I__11617\ : InMux
    port map (
            O => \N__50662\,
            I => \N__50654\
        );

    \I__11616\ : Span4Mux_h
    port map (
            O => \N__50657\,
            I => \N__50651\
        );

    \I__11615\ : LocalMux
    port map (
            O => \N__50654\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__11614\ : Odrv4
    port map (
            O => \N__50651\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__11613\ : InMux
    port map (
            O => \N__50646\,
            I => \N__50643\
        );

    \I__11612\ : LocalMux
    port map (
            O => \N__50643\,
            I => \N__50640\
        );

    \I__11611\ : Span4Mux_h
    port map (
            O => \N__50640\,
            I => \N__50636\
        );

    \I__11610\ : InMux
    port map (
            O => \N__50639\,
            I => \N__50633\
        );

    \I__11609\ : Odrv4
    port map (
            O => \N__50636\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__11608\ : LocalMux
    port map (
            O => \N__50633\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__11607\ : CascadeMux
    port map (
            O => \N__50628\,
            I => \N__50624\
        );

    \I__11606\ : InMux
    port map (
            O => \N__50627\,
            I => \N__50621\
        );

    \I__11605\ : InMux
    port map (
            O => \N__50624\,
            I => \N__50618\
        );

    \I__11604\ : LocalMux
    port map (
            O => \N__50621\,
            I => \N__50612\
        );

    \I__11603\ : LocalMux
    port map (
            O => \N__50618\,
            I => \N__50612\
        );

    \I__11602\ : InMux
    port map (
            O => \N__50617\,
            I => \N__50609\
        );

    \I__11601\ : Span4Mux_h
    port map (
            O => \N__50612\,
            I => \N__50606\
        );

    \I__11600\ : LocalMux
    port map (
            O => \N__50609\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__11599\ : Odrv4
    port map (
            O => \N__50606\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__11598\ : InMux
    port map (
            O => \N__50601\,
            I => \N__50598\
        );

    \I__11597\ : LocalMux
    port map (
            O => \N__50598\,
            I => \N__50595\
        );

    \I__11596\ : Span4Mux_v
    port map (
            O => \N__50595\,
            I => \N__50591\
        );

    \I__11595\ : InMux
    port map (
            O => \N__50594\,
            I => \N__50588\
        );

    \I__11594\ : Odrv4
    port map (
            O => \N__50591\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__50588\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__11592\ : CEMux
    port map (
            O => \N__50583\,
            I => \N__50579\
        );

    \I__11591\ : CEMux
    port map (
            O => \N__50582\,
            I => \N__50576\
        );

    \I__11590\ : LocalMux
    port map (
            O => \N__50579\,
            I => \N__50570\
        );

    \I__11589\ : LocalMux
    port map (
            O => \N__50576\,
            I => \N__50567\
        );

    \I__11588\ : CEMux
    port map (
            O => \N__50575\,
            I => \N__50564\
        );

    \I__11587\ : CEMux
    port map (
            O => \N__50574\,
            I => \N__50561\
        );

    \I__11586\ : CEMux
    port map (
            O => \N__50573\,
            I => \N__50558\
        );

    \I__11585\ : Span4Mux_h
    port map (
            O => \N__50570\,
            I => \N__50549\
        );

    \I__11584\ : Span4Mux_v
    port map (
            O => \N__50567\,
            I => \N__50549\
        );

    \I__11583\ : LocalMux
    port map (
            O => \N__50564\,
            I => \N__50549\
        );

    \I__11582\ : LocalMux
    port map (
            O => \N__50561\,
            I => \N__50549\
        );

    \I__11581\ : LocalMux
    port map (
            O => \N__50558\,
            I => \N__50546\
        );

    \I__11580\ : Odrv4
    port map (
            O => \N__50549\,
            I => \delay_measurement_inst.delay_hc_timer.N_155_i\
        );

    \I__11579\ : Odrv4
    port map (
            O => \N__50546\,
            I => \delay_measurement_inst.delay_hc_timer.N_155_i\
        );

    \I__11578\ : InMux
    port map (
            O => \N__50541\,
            I => \N__50538\
        );

    \I__11577\ : LocalMux
    port map (
            O => \N__50538\,
            I => \N__50535\
        );

    \I__11576\ : Span4Mux_v
    port map (
            O => \N__50535\,
            I => \N__50532\
        );

    \I__11575\ : Span4Mux_h
    port map (
            O => \N__50532\,
            I => \N__50529\
        );

    \I__11574\ : Odrv4
    port map (
            O => \N__50529\,
            I => \pwm_generator_inst.O_0\
        );

    \I__11573\ : InMux
    port map (
            O => \N__50526\,
            I => \N__50523\
        );

    \I__11572\ : LocalMux
    port map (
            O => \N__50523\,
            I => \pwm_generator_inst.un15_threshold_1_axb_0\
        );

    \I__11571\ : InMux
    port map (
            O => \N__50520\,
            I => \N__50517\
        );

    \I__11570\ : LocalMux
    port map (
            O => \N__50517\,
            I => \N__50514\
        );

    \I__11569\ : Span12Mux_s7_v
    port map (
            O => \N__50514\,
            I => \N__50511\
        );

    \I__11568\ : Odrv12
    port map (
            O => \N__50511\,
            I => \pwm_generator_inst.O_1\
        );

    \I__11567\ : InMux
    port map (
            O => \N__50508\,
            I => \N__50505\
        );

    \I__11566\ : LocalMux
    port map (
            O => \N__50505\,
            I => \pwm_generator_inst.un15_threshold_1_axb_1\
        );

    \I__11565\ : InMux
    port map (
            O => \N__50502\,
            I => \N__50499\
        );

    \I__11564\ : LocalMux
    port map (
            O => \N__50499\,
            I => \N__50496\
        );

    \I__11563\ : Span12Mux_h
    port map (
            O => \N__50496\,
            I => \N__50493\
        );

    \I__11562\ : Odrv12
    port map (
            O => \N__50493\,
            I => \pwm_generator_inst.O_2\
        );

    \I__11561\ : InMux
    port map (
            O => \N__50490\,
            I => \N__50487\
        );

    \I__11560\ : LocalMux
    port map (
            O => \N__50487\,
            I => \pwm_generator_inst.un15_threshold_1_axb_2\
        );

    \I__11559\ : InMux
    port map (
            O => \N__50484\,
            I => \N__50481\
        );

    \I__11558\ : LocalMux
    port map (
            O => \N__50481\,
            I => \N__50478\
        );

    \I__11557\ : Span4Mux_v
    port map (
            O => \N__50478\,
            I => \N__50474\
        );

    \I__11556\ : InMux
    port map (
            O => \N__50477\,
            I => \N__50471\
        );

    \I__11555\ : Odrv4
    port map (
            O => \N__50474\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__50471\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__11553\ : InMux
    port map (
            O => \N__50466\,
            I => \N__50463\
        );

    \I__11552\ : LocalMux
    port map (
            O => \N__50463\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__11551\ : CascadeMux
    port map (
            O => \N__50460\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\
        );

    \I__11550\ : InMux
    port map (
            O => \N__50457\,
            I => \N__50454\
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__50454\,
            I => \N__50451\
        );

    \I__11548\ : Odrv4
    port map (
            O => \N__50451\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23\
        );

    \I__11547\ : InMux
    port map (
            O => \N__50448\,
            I => \N__50444\
        );

    \I__11546\ : InMux
    port map (
            O => \N__50447\,
            I => \N__50441\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__50444\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__50441\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__11543\ : InMux
    port map (
            O => \N__50436\,
            I => \N__50433\
        );

    \I__11542\ : LocalMux
    port map (
            O => \N__50433\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13\
        );

    \I__11541\ : InMux
    port map (
            O => \N__50430\,
            I => \N__50427\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__50427\,
            I => \N__50423\
        );

    \I__11539\ : InMux
    port map (
            O => \N__50426\,
            I => \N__50420\
        );

    \I__11538\ : Odrv4
    port map (
            O => \N__50423\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__11537\ : LocalMux
    port map (
            O => \N__50420\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__11536\ : InMux
    port map (
            O => \N__50415\,
            I => \N__50411\
        );

    \I__11535\ : InMux
    port map (
            O => \N__50414\,
            I => \N__50408\
        );

    \I__11534\ : LocalMux
    port map (
            O => \N__50411\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__11533\ : LocalMux
    port map (
            O => \N__50408\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__11532\ : InMux
    port map (
            O => \N__50403\,
            I => \N__50400\
        );

    \I__11531\ : LocalMux
    port map (
            O => \N__50400\,
            I => \N__50397\
        );

    \I__11530\ : Span4Mux_v
    port map (
            O => \N__50397\,
            I => \N__50393\
        );

    \I__11529\ : InMux
    port map (
            O => \N__50396\,
            I => \N__50390\
        );

    \I__11528\ : Odrv4
    port map (
            O => \N__50393\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__11527\ : LocalMux
    port map (
            O => \N__50390\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__11526\ : InMux
    port map (
            O => \N__50385\,
            I => \N__50382\
        );

    \I__11525\ : LocalMux
    port map (
            O => \N__50382\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__11524\ : CascadeMux
    port map (
            O => \N__50379\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27_cascade_\
        );

    \I__11523\ : InMux
    port map (
            O => \N__50376\,
            I => \N__50373\
        );

    \I__11522\ : LocalMux
    port map (
            O => \N__50373\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27\
        );

    \I__11521\ : InMux
    port map (
            O => \N__50370\,
            I => \N__50366\
        );

    \I__11520\ : InMux
    port map (
            O => \N__50369\,
            I => \N__50363\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__50366\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__11518\ : LocalMux
    port map (
            O => \N__50363\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__11517\ : InMux
    port map (
            O => \N__50358\,
            I => \N__50355\
        );

    \I__11516\ : LocalMux
    port map (
            O => \N__50355\,
            I => \N__50351\
        );

    \I__11515\ : InMux
    port map (
            O => \N__50354\,
            I => \N__50348\
        );

    \I__11514\ : Odrv4
    port map (
            O => \N__50351\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__11513\ : LocalMux
    port map (
            O => \N__50348\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__11512\ : InMux
    port map (
            O => \N__50343\,
            I => \N__50340\
        );

    \I__11511\ : LocalMux
    port map (
            O => \N__50340\,
            I => \N__50337\
        );

    \I__11510\ : Span4Mux_h
    port map (
            O => \N__50337\,
            I => \N__50333\
        );

    \I__11509\ : InMux
    port map (
            O => \N__50336\,
            I => \N__50330\
        );

    \I__11508\ : Odrv4
    port map (
            O => \N__50333\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__50330\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__11506\ : InMux
    port map (
            O => \N__50325\,
            I => \N__50322\
        );

    \I__11505\ : LocalMux
    port map (
            O => \N__50322\,
            I => \N__50318\
        );

    \I__11504\ : InMux
    port map (
            O => \N__50321\,
            I => \N__50315\
        );

    \I__11503\ : Odrv4
    port map (
            O => \N__50318\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__50315\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__11501\ : CascadeMux
    port map (
            O => \N__50310\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_\
        );

    \I__11500\ : InMux
    port map (
            O => \N__50307\,
            I => \N__50300\
        );

    \I__11499\ : InMux
    port map (
            O => \N__50306\,
            I => \N__50300\
        );

    \I__11498\ : InMux
    port map (
            O => \N__50305\,
            I => \N__50297\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__50300\,
            I => \N__50294\
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__50297\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_26\
        );

    \I__11495\ : Odrv12
    port map (
            O => \N__50294\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_26\
        );

    \I__11494\ : CascadeMux
    port map (
            O => \N__50289\,
            I => \N__50285\
        );

    \I__11493\ : CascadeMux
    port map (
            O => \N__50288\,
            I => \N__50282\
        );

    \I__11492\ : InMux
    port map (
            O => \N__50285\,
            I => \N__50277\
        );

    \I__11491\ : InMux
    port map (
            O => \N__50282\,
            I => \N__50277\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__50277\,
            I => \N__50273\
        );

    \I__11489\ : InMux
    port map (
            O => \N__50276\,
            I => \N__50270\
        );

    \I__11488\ : Span4Mux_h
    port map (
            O => \N__50273\,
            I => \N__50267\
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__50270\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_27\
        );

    \I__11486\ : Odrv4
    port map (
            O => \N__50267\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_27\
        );

    \I__11485\ : CascadeMux
    port map (
            O => \N__50262\,
            I => \N__50259\
        );

    \I__11484\ : InMux
    port map (
            O => \N__50259\,
            I => \N__50256\
        );

    \I__11483\ : LocalMux
    port map (
            O => \N__50256\,
            I => \N__50253\
        );

    \I__11482\ : Span4Mux_h
    port map (
            O => \N__50253\,
            I => \N__50250\
        );

    \I__11481\ : Odrv4
    port map (
            O => \N__50250\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26\
        );

    \I__11480\ : InMux
    port map (
            O => \N__50247\,
            I => \N__50243\
        );

    \I__11479\ : InMux
    port map (
            O => \N__50246\,
            I => \N__50240\
        );

    \I__11478\ : LocalMux
    port map (
            O => \N__50243\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_27
        );

    \I__11477\ : LocalMux
    port map (
            O => \N__50240\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_27
        );

    \I__11476\ : InMux
    port map (
            O => \N__50235\,
            I => \N__50229\
        );

    \I__11475\ : InMux
    port map (
            O => \N__50234\,
            I => \N__50229\
        );

    \I__11474\ : LocalMux
    port map (
            O => \N__50229\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_27\
        );

    \I__11473\ : InMux
    port map (
            O => \N__50226\,
            I => \N__50222\
        );

    \I__11472\ : InMux
    port map (
            O => \N__50225\,
            I => \N__50219\
        );

    \I__11471\ : LocalMux
    port map (
            O => \N__50222\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_26
        );

    \I__11470\ : LocalMux
    port map (
            O => \N__50219\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_26
        );

    \I__11469\ : InMux
    port map (
            O => \N__50214\,
            I => \N__50208\
        );

    \I__11468\ : InMux
    port map (
            O => \N__50213\,
            I => \N__50208\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__50208\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_26\
        );

    \I__11466\ : InMux
    port map (
            O => \N__50205\,
            I => \N__50201\
        );

    \I__11465\ : InMux
    port map (
            O => \N__50204\,
            I => \N__50198\
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__50201\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_24
        );

    \I__11463\ : LocalMux
    port map (
            O => \N__50198\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_24
        );

    \I__11462\ : InMux
    port map (
            O => \N__50193\,
            I => \N__50187\
        );

    \I__11461\ : InMux
    port map (
            O => \N__50192\,
            I => \N__50187\
        );

    \I__11460\ : LocalMux
    port map (
            O => \N__50187\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_24\
        );

    \I__11459\ : InMux
    port map (
            O => \N__50184\,
            I => \N__50180\
        );

    \I__11458\ : InMux
    port map (
            O => \N__50183\,
            I => \N__50177\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__50180\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_25
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__50177\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_25
        );

    \I__11455\ : CascadeMux
    port map (
            O => \N__50172\,
            I => \N__50168\
        );

    \I__11454\ : CascadeMux
    port map (
            O => \N__50171\,
            I => \N__50165\
        );

    \I__11453\ : InMux
    port map (
            O => \N__50168\,
            I => \N__50160\
        );

    \I__11452\ : InMux
    port map (
            O => \N__50165\,
            I => \N__50160\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__50160\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_25\
        );

    \I__11450\ : CEMux
    port map (
            O => \N__50157\,
            I => \N__50152\
        );

    \I__11449\ : CEMux
    port map (
            O => \N__50156\,
            I => \N__50149\
        );

    \I__11448\ : CEMux
    port map (
            O => \N__50155\,
            I => \N__50142\
        );

    \I__11447\ : LocalMux
    port map (
            O => \N__50152\,
            I => \N__50135\
        );

    \I__11446\ : LocalMux
    port map (
            O => \N__50149\,
            I => \N__50135\
        );

    \I__11445\ : CEMux
    port map (
            O => \N__50148\,
            I => \N__50132\
        );

    \I__11444\ : CEMux
    port map (
            O => \N__50147\,
            I => \N__50128\
        );

    \I__11443\ : CEMux
    port map (
            O => \N__50146\,
            I => \N__50125\
        );

    \I__11442\ : CEMux
    port map (
            O => \N__50145\,
            I => \N__50122\
        );

    \I__11441\ : LocalMux
    port map (
            O => \N__50142\,
            I => \N__50119\
        );

    \I__11440\ : CEMux
    port map (
            O => \N__50141\,
            I => \N__50116\
        );

    \I__11439\ : CEMux
    port map (
            O => \N__50140\,
            I => \N__50113\
        );

    \I__11438\ : Span4Mux_v
    port map (
            O => \N__50135\,
            I => \N__50108\
        );

    \I__11437\ : LocalMux
    port map (
            O => \N__50132\,
            I => \N__50108\
        );

    \I__11436\ : CEMux
    port map (
            O => \N__50131\,
            I => \N__50105\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__50128\,
            I => \N__50098\
        );

    \I__11434\ : LocalMux
    port map (
            O => \N__50125\,
            I => \N__50098\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__50122\,
            I => \N__50098\
        );

    \I__11432\ : Span4Mux_v
    port map (
            O => \N__50119\,
            I => \N__50095\
        );

    \I__11431\ : LocalMux
    port map (
            O => \N__50116\,
            I => \N__50088\
        );

    \I__11430\ : LocalMux
    port map (
            O => \N__50113\,
            I => \N__50088\
        );

    \I__11429\ : Span4Mux_v
    port map (
            O => \N__50108\,
            I => \N__50088\
        );

    \I__11428\ : LocalMux
    port map (
            O => \N__50105\,
            I => \N__50085\
        );

    \I__11427\ : Span4Mux_v
    port map (
            O => \N__50098\,
            I => \N__50082\
        );

    \I__11426\ : Span4Mux_v
    port map (
            O => \N__50095\,
            I => \N__50077\
        );

    \I__11425\ : Span4Mux_v
    port map (
            O => \N__50088\,
            I => \N__50077\
        );

    \I__11424\ : Span12Mux_v
    port map (
            O => \N__50085\,
            I => \N__50074\
        );

    \I__11423\ : Span4Mux_h
    port map (
            O => \N__50082\,
            I => \N__50071\
        );

    \I__11422\ : Span4Mux_h
    port map (
            O => \N__50077\,
            I => \N__50068\
        );

    \I__11421\ : Odrv12
    port map (
            O => \N__50074\,
            I => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__11420\ : Odrv4
    port map (
            O => \N__50071\,
            I => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__11419\ : Odrv4
    port map (
            O => \N__50068\,
            I => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__11418\ : InMux
    port map (
            O => \N__50061\,
            I => \N__50058\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__50058\,
            I => \N__50054\
        );

    \I__11416\ : CascadeMux
    port map (
            O => \N__50057\,
            I => \N__50051\
        );

    \I__11415\ : Span4Mux_v
    port map (
            O => \N__50054\,
            I => \N__50048\
        );

    \I__11414\ : InMux
    port map (
            O => \N__50051\,
            I => \N__50045\
        );

    \I__11413\ : Odrv4
    port map (
            O => \N__50048\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__11412\ : LocalMux
    port map (
            O => \N__50045\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__11411\ : InMux
    port map (
            O => \N__50040\,
            I => \N__50037\
        );

    \I__11410\ : LocalMux
    port map (
            O => \N__50037\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__11409\ : CascadeMux
    port map (
            O => \N__50034\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12_cascade_\
        );

    \I__11408\ : InMux
    port map (
            O => \N__50031\,
            I => \N__50028\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__50028\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12\
        );

    \I__11406\ : InMux
    port map (
            O => \N__50025\,
            I => \N__50022\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__50022\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5\
        );

    \I__11404\ : InMux
    port map (
            O => \N__50019\,
            I => \N__50016\
        );

    \I__11403\ : LocalMux
    port map (
            O => \N__50016\,
            I => \N__50012\
        );

    \I__11402\ : InMux
    port map (
            O => \N__50015\,
            I => \N__50009\
        );

    \I__11401\ : Odrv4
    port map (
            O => \N__50012\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_19
        );

    \I__11400\ : LocalMux
    port map (
            O => \N__50009\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_19
        );

    \I__11399\ : InMux
    port map (
            O => \N__50004\,
            I => \N__50001\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__50001\,
            I => \N__49998\
        );

    \I__11397\ : Span4Mux_h
    port map (
            O => \N__49998\,
            I => \N__49995\
        );

    \I__11396\ : Odrv4
    port map (
            O => \N__49995\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt16\
        );

    \I__11395\ : InMux
    port map (
            O => \N__49992\,
            I => \N__49986\
        );

    \I__11394\ : InMux
    port map (
            O => \N__49991\,
            I => \N__49986\
        );

    \I__11393\ : LocalMux
    port map (
            O => \N__49986\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_16\
        );

    \I__11392\ : InMux
    port map (
            O => \N__49983\,
            I => \N__49976\
        );

    \I__11391\ : InMux
    port map (
            O => \N__49982\,
            I => \N__49976\
        );

    \I__11390\ : InMux
    port map (
            O => \N__49981\,
            I => \N__49973\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__49976\,
            I => \N__49970\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__49973\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_17\
        );

    \I__11387\ : Odrv12
    port map (
            O => \N__49970\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_17\
        );

    \I__11386\ : CascadeMux
    port map (
            O => \N__49965\,
            I => \N__49961\
        );

    \I__11385\ : CascadeMux
    port map (
            O => \N__49964\,
            I => \N__49958\
        );

    \I__11384\ : InMux
    port map (
            O => \N__49961\,
            I => \N__49952\
        );

    \I__11383\ : InMux
    port map (
            O => \N__49958\,
            I => \N__49952\
        );

    \I__11382\ : InMux
    port map (
            O => \N__49957\,
            I => \N__49949\
        );

    \I__11381\ : LocalMux
    port map (
            O => \N__49952\,
            I => \N__49946\
        );

    \I__11380\ : LocalMux
    port map (
            O => \N__49949\,
            I => \N__49941\
        );

    \I__11379\ : Span4Mux_h
    port map (
            O => \N__49946\,
            I => \N__49941\
        );

    \I__11378\ : Odrv4
    port map (
            O => \N__49941\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_16\
        );

    \I__11377\ : CascadeMux
    port map (
            O => \N__49938\,
            I => \N__49935\
        );

    \I__11376\ : InMux
    port map (
            O => \N__49935\,
            I => \N__49932\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__49932\,
            I => \N__49929\
        );

    \I__11374\ : Span4Mux_h
    port map (
            O => \N__49929\,
            I => \N__49926\
        );

    \I__11373\ : Odrv4
    port map (
            O => \N__49926\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16\
        );

    \I__11372\ : InMux
    port map (
            O => \N__49923\,
            I => \N__49920\
        );

    \I__11371\ : LocalMux
    port map (
            O => \N__49920\,
            I => \N__49917\
        );

    \I__11370\ : Span4Mux_v
    port map (
            O => \N__49917\,
            I => \N__49913\
        );

    \I__11369\ : InMux
    port map (
            O => \N__49916\,
            I => \N__49910\
        );

    \I__11368\ : Odrv4
    port map (
            O => \N__49913\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_17
        );

    \I__11367\ : LocalMux
    port map (
            O => \N__49910\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_17
        );

    \I__11366\ : InMux
    port map (
            O => \N__49905\,
            I => \N__49899\
        );

    \I__11365\ : InMux
    port map (
            O => \N__49904\,
            I => \N__49899\
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__49899\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_17\
        );

    \I__11363\ : CascadeMux
    port map (
            O => \N__49896\,
            I => \N__49893\
        );

    \I__11362\ : InMux
    port map (
            O => \N__49893\,
            I => \N__49890\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__49890\,
            I => \N__49887\
        );

    \I__11360\ : Span4Mux_v
    port map (
            O => \N__49887\,
            I => \N__49884\
        );

    \I__11359\ : Odrv4
    port map (
            O => \N__49884\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt18\
        );

    \I__11358\ : InMux
    port map (
            O => \N__49881\,
            I => \N__49875\
        );

    \I__11357\ : InMux
    port map (
            O => \N__49880\,
            I => \N__49875\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__49875\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18\
        );

    \I__11355\ : InMux
    port map (
            O => \N__49872\,
            I => \N__49866\
        );

    \I__11354\ : InMux
    port map (
            O => \N__49871\,
            I => \N__49866\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__49866\,
            I => \N__49862\
        );

    \I__11352\ : InMux
    port map (
            O => \N__49865\,
            I => \N__49859\
        );

    \I__11351\ : Span4Mux_h
    port map (
            O => \N__49862\,
            I => \N__49856\
        );

    \I__11350\ : LocalMux
    port map (
            O => \N__49859\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_19\
        );

    \I__11349\ : Odrv4
    port map (
            O => \N__49856\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_19\
        );

    \I__11348\ : CascadeMux
    port map (
            O => \N__49851\,
            I => \N__49847\
        );

    \I__11347\ : CascadeMux
    port map (
            O => \N__49850\,
            I => \N__49844\
        );

    \I__11346\ : InMux
    port map (
            O => \N__49847\,
            I => \N__49838\
        );

    \I__11345\ : InMux
    port map (
            O => \N__49844\,
            I => \N__49838\
        );

    \I__11344\ : InMux
    port map (
            O => \N__49843\,
            I => \N__49835\
        );

    \I__11343\ : LocalMux
    port map (
            O => \N__49838\,
            I => \N__49832\
        );

    \I__11342\ : LocalMux
    port map (
            O => \N__49835\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_18\
        );

    \I__11341\ : Odrv12
    port map (
            O => \N__49832\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_18\
        );

    \I__11340\ : InMux
    port map (
            O => \N__49827\,
            I => \N__49821\
        );

    \I__11339\ : InMux
    port map (
            O => \N__49826\,
            I => \N__49821\
        );

    \I__11338\ : LocalMux
    port map (
            O => \N__49821\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19\
        );

    \I__11337\ : InMux
    port map (
            O => \N__49818\,
            I => \N__49815\
        );

    \I__11336\ : LocalMux
    port map (
            O => \N__49815\,
            I => \N__49812\
        );

    \I__11335\ : Span4Mux_h
    port map (
            O => \N__49812\,
            I => \N__49809\
        );

    \I__11334\ : Odrv4
    port map (
            O => \N__49809\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18\
        );

    \I__11333\ : CascadeMux
    port map (
            O => \N__49806\,
            I => \N__49803\
        );

    \I__11332\ : InMux
    port map (
            O => \N__49803\,
            I => \N__49800\
        );

    \I__11331\ : LocalMux
    port map (
            O => \N__49800\,
            I => \N__49797\
        );

    \I__11330\ : Span4Mux_h
    port map (
            O => \N__49797\,
            I => \N__49794\
        );

    \I__11329\ : Odrv4
    port map (
            O => \N__49794\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt24\
        );

    \I__11328\ : InMux
    port map (
            O => \N__49791\,
            I => \N__49784\
        );

    \I__11327\ : InMux
    port map (
            O => \N__49790\,
            I => \N__49784\
        );

    \I__11326\ : InMux
    port map (
            O => \N__49789\,
            I => \N__49781\
        );

    \I__11325\ : LocalMux
    port map (
            O => \N__49784\,
            I => \N__49778\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__49781\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_25\
        );

    \I__11323\ : Odrv12
    port map (
            O => \N__49778\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_25\
        );

    \I__11322\ : InMux
    port map (
            O => \N__49773\,
            I => \N__49766\
        );

    \I__11321\ : InMux
    port map (
            O => \N__49772\,
            I => \N__49766\
        );

    \I__11320\ : InMux
    port map (
            O => \N__49771\,
            I => \N__49763\
        );

    \I__11319\ : LocalMux
    port map (
            O => \N__49766\,
            I => \N__49760\
        );

    \I__11318\ : LocalMux
    port map (
            O => \N__49763\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_24\
        );

    \I__11317\ : Odrv12
    port map (
            O => \N__49760\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_24\
        );

    \I__11316\ : InMux
    port map (
            O => \N__49755\,
            I => \N__49752\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__49752\,
            I => \N__49749\
        );

    \I__11314\ : Odrv12
    port map (
            O => \N__49749\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24\
        );

    \I__11313\ : InMux
    port map (
            O => \N__49746\,
            I => \N__49743\
        );

    \I__11312\ : LocalMux
    port map (
            O => \N__49743\,
            I => \N__49740\
        );

    \I__11311\ : Odrv12
    port map (
            O => \N__49740\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt26\
        );

    \I__11310\ : InMux
    port map (
            O => \N__49737\,
            I => \N__49734\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__49734\,
            I => \pwm_generator_inst.un19_threshold_0_axb_7\
        );

    \I__11308\ : CascadeMux
    port map (
            O => \N__49731\,
            I => \N__49728\
        );

    \I__11307\ : InMux
    port map (
            O => \N__49728\,
            I => \N__49725\
        );

    \I__11306\ : LocalMux
    port map (
            O => \N__49725\,
            I => \N__49722\
        );

    \I__11305\ : Span4Mux_v
    port map (
            O => \N__49722\,
            I => \N__49719\
        );

    \I__11304\ : Odrv4
    port map (
            O => \N__49719\,
            I => \pwm_generator_inst.un14_counter_7\
        );

    \I__11303\ : InMux
    port map (
            O => \N__49716\,
            I => \pwm_generator_inst.un19_threshold_0_cry_6\
        );

    \I__11302\ : CascadeMux
    port map (
            O => \N__49713\,
            I => \N__49710\
        );

    \I__11301\ : InMux
    port map (
            O => \N__49710\,
            I => \N__49707\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__49707\,
            I => \N__49704\
        );

    \I__11299\ : Odrv12
    port map (
            O => \N__49704\,
            I => \pwm_generator_inst.un14_counter_8\
        );

    \I__11298\ : InMux
    port map (
            O => \N__49701\,
            I => \bfn_17_27_0_\
        );

    \I__11297\ : InMux
    port map (
            O => \N__49698\,
            I => \N__49695\
        );

    \I__11296\ : LocalMux
    port map (
            O => \N__49695\,
            I => \N__49692\
        );

    \I__11295\ : Span4Mux_h
    port map (
            O => \N__49692\,
            I => \N__49689\
        );

    \I__11294\ : Odrv4
    port map (
            O => \N__49689\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\
        );

    \I__11293\ : InMux
    port map (
            O => \N__49686\,
            I => \pwm_generator_inst.un19_threshold_0_cry_8\
        );

    \I__11292\ : CascadeMux
    port map (
            O => \N__49683\,
            I => \N__49680\
        );

    \I__11291\ : InMux
    port map (
            O => \N__49680\,
            I => \N__49677\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__49677\,
            I => \N__49674\
        );

    \I__11289\ : Odrv4
    port map (
            O => \N__49674\,
            I => \pwm_generator_inst.un14_counter_9\
        );

    \I__11288\ : InMux
    port map (
            O => \N__49671\,
            I => \N__49668\
        );

    \I__11287\ : LocalMux
    port map (
            O => \N__49668\,
            I => \N__49665\
        );

    \I__11286\ : Span4Mux_h
    port map (
            O => \N__49665\,
            I => \N__49661\
        );

    \I__11285\ : InMux
    port map (
            O => \N__49664\,
            I => \N__49658\
        );

    \I__11284\ : Odrv4
    port map (
            O => \N__49661\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__11283\ : LocalMux
    port map (
            O => \N__49658\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__11282\ : InMux
    port map (
            O => \N__49653\,
            I => \N__49650\
        );

    \I__11281\ : LocalMux
    port map (
            O => \N__49650\,
            I => \pwm_generator_inst.un19_threshold_0_axb_6\
        );

    \I__11280\ : CascadeMux
    port map (
            O => \N__49647\,
            I => \N__49644\
        );

    \I__11279\ : InMux
    port map (
            O => \N__49644\,
            I => \N__49641\
        );

    \I__11278\ : LocalMux
    port map (
            O => \N__49641\,
            I => \N__49637\
        );

    \I__11277\ : InMux
    port map (
            O => \N__49640\,
            I => \N__49634\
        );

    \I__11276\ : Span4Mux_h
    port map (
            O => \N__49637\,
            I => \N__49631\
        );

    \I__11275\ : LocalMux
    port map (
            O => \N__49634\,
            I => \N__49628\
        );

    \I__11274\ : Odrv4
    port map (
            O => \N__49631\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__11273\ : Odrv4
    port map (
            O => \N__49628\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__11272\ : InMux
    port map (
            O => \N__49623\,
            I => \N__49620\
        );

    \I__11271\ : LocalMux
    port map (
            O => \N__49620\,
            I => \pwm_generator_inst.un19_threshold_0_axb_4\
        );

    \I__11270\ : InMux
    port map (
            O => \N__49617\,
            I => \N__49614\
        );

    \I__11269\ : LocalMux
    port map (
            O => \N__49614\,
            I => \N__49611\
        );

    \I__11268\ : Span4Mux_h
    port map (
            O => \N__49611\,
            I => \N__49607\
        );

    \I__11267\ : InMux
    port map (
            O => \N__49610\,
            I => \N__49604\
        );

    \I__11266\ : Odrv4
    port map (
            O => \N__49607\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__11265\ : LocalMux
    port map (
            O => \N__49604\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__11264\ : InMux
    port map (
            O => \N__49599\,
            I => \N__49596\
        );

    \I__11263\ : LocalMux
    port map (
            O => \N__49596\,
            I => \pwm_generator_inst.un19_threshold_0_axb_8\
        );

    \I__11262\ : InMux
    port map (
            O => \N__49593\,
            I => \N__49590\
        );

    \I__11261\ : LocalMux
    port map (
            O => \N__49590\,
            I => \N__49586\
        );

    \I__11260\ : InMux
    port map (
            O => \N__49589\,
            I => \N__49583\
        );

    \I__11259\ : Odrv4
    port map (
            O => \N__49586\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_16
        );

    \I__11258\ : LocalMux
    port map (
            O => \N__49583\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_16
        );

    \I__11257\ : InMux
    port map (
            O => \N__49578\,
            I => \N__49574\
        );

    \I__11256\ : InMux
    port map (
            O => \N__49577\,
            I => \N__49571\
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__49574\,
            I => \N__49568\
        );

    \I__11254\ : LocalMux
    port map (
            O => \N__49571\,
            I => \N__49565\
        );

    \I__11253\ : Span4Mux_h
    port map (
            O => \N__49568\,
            I => \N__49562\
        );

    \I__11252\ : Odrv4
    port map (
            O => \N__49565\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_18
        );

    \I__11251\ : Odrv4
    port map (
            O => \N__49562\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_18
        );

    \I__11250\ : InMux
    port map (
            O => \N__49557\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__11249\ : IoInMux
    port map (
            O => \N__49554\,
            I => \N__49551\
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__49551\,
            I => \N__49548\
        );

    \I__11247\ : Span4Mux_s0_v
    port map (
            O => \N__49548\,
            I => \N__49545\
        );

    \I__11246\ : Sp12to4
    port map (
            O => \N__49545\,
            I => \N__49542\
        );

    \I__11245\ : Span12Mux_h
    port map (
            O => \N__49542\,
            I => \N__49539\
        );

    \I__11244\ : Span12Mux_v
    port map (
            O => \N__49539\,
            I => \N__49536\
        );

    \I__11243\ : Span12Mux_v
    port map (
            O => \N__49536\,
            I => \N__49533\
        );

    \I__11242\ : Odrv12
    port map (
            O => \N__49533\,
            I => pwm_output_c
        );

    \I__11241\ : InMux
    port map (
            O => \N__49530\,
            I => \N__49527\
        );

    \I__11240\ : LocalMux
    port map (
            O => \N__49527\,
            I => \pwm_generator_inst.un19_threshold_0_axb_0\
        );

    \I__11239\ : CascadeMux
    port map (
            O => \N__49524\,
            I => \N__49521\
        );

    \I__11238\ : InMux
    port map (
            O => \N__49521\,
            I => \N__49518\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__49518\,
            I => \N__49515\
        );

    \I__11236\ : Span4Mux_h
    port map (
            O => \N__49515\,
            I => \N__49512\
        );

    \I__11235\ : Odrv4
    port map (
            O => \N__49512\,
            I => \pwm_generator_inst.un14_counter_0\
        );

    \I__11234\ : CascadeMux
    port map (
            O => \N__49509\,
            I => \N__49506\
        );

    \I__11233\ : InMux
    port map (
            O => \N__49506\,
            I => \N__49503\
        );

    \I__11232\ : LocalMux
    port map (
            O => \N__49503\,
            I => \N__49500\
        );

    \I__11231\ : Span4Mux_h
    port map (
            O => \N__49500\,
            I => \N__49497\
        );

    \I__11230\ : Odrv4
    port map (
            O => \N__49497\,
            I => \pwm_generator_inst.un14_counter_1\
        );

    \I__11229\ : InMux
    port map (
            O => \N__49494\,
            I => \pwm_generator_inst.un19_threshold_0_cry_0\
        );

    \I__11228\ : CascadeMux
    port map (
            O => \N__49491\,
            I => \N__49488\
        );

    \I__11227\ : InMux
    port map (
            O => \N__49488\,
            I => \N__49485\
        );

    \I__11226\ : LocalMux
    port map (
            O => \N__49485\,
            I => \pwm_generator_inst.un19_threshold_0_axb_2\
        );

    \I__11225\ : CascadeMux
    port map (
            O => \N__49482\,
            I => \N__49479\
        );

    \I__11224\ : InMux
    port map (
            O => \N__49479\,
            I => \N__49476\
        );

    \I__11223\ : LocalMux
    port map (
            O => \N__49476\,
            I => \N__49473\
        );

    \I__11222\ : Span4Mux_v
    port map (
            O => \N__49473\,
            I => \N__49470\
        );

    \I__11221\ : Odrv4
    port map (
            O => \N__49470\,
            I => \pwm_generator_inst.un14_counter_2\
        );

    \I__11220\ : InMux
    port map (
            O => \N__49467\,
            I => \pwm_generator_inst.un19_threshold_0_cry_1\
        );

    \I__11219\ : InMux
    port map (
            O => \N__49464\,
            I => \N__49461\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__49461\,
            I => \pwm_generator_inst.un19_threshold_0_axb_3\
        );

    \I__11217\ : CascadeMux
    port map (
            O => \N__49458\,
            I => \N__49455\
        );

    \I__11216\ : InMux
    port map (
            O => \N__49455\,
            I => \N__49452\
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__49452\,
            I => \N__49449\
        );

    \I__11214\ : Span4Mux_v
    port map (
            O => \N__49449\,
            I => \N__49446\
        );

    \I__11213\ : Odrv4
    port map (
            O => \N__49446\,
            I => \pwm_generator_inst.un14_counter_3\
        );

    \I__11212\ : InMux
    port map (
            O => \N__49443\,
            I => \pwm_generator_inst.un19_threshold_0_cry_2\
        );

    \I__11211\ : CascadeMux
    port map (
            O => \N__49440\,
            I => \N__49437\
        );

    \I__11210\ : InMux
    port map (
            O => \N__49437\,
            I => \N__49434\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__49434\,
            I => \N__49431\
        );

    \I__11208\ : Odrv4
    port map (
            O => \N__49431\,
            I => \pwm_generator_inst.un14_counter_4\
        );

    \I__11207\ : InMux
    port map (
            O => \N__49428\,
            I => \pwm_generator_inst.un19_threshold_0_cry_3\
        );

    \I__11206\ : InMux
    port map (
            O => \N__49425\,
            I => \N__49422\
        );

    \I__11205\ : LocalMux
    port map (
            O => \N__49422\,
            I => \pwm_generator_inst.un19_threshold_0_axb_5\
        );

    \I__11204\ : CascadeMux
    port map (
            O => \N__49419\,
            I => \N__49416\
        );

    \I__11203\ : InMux
    port map (
            O => \N__49416\,
            I => \N__49413\
        );

    \I__11202\ : LocalMux
    port map (
            O => \N__49413\,
            I => \N__49410\
        );

    \I__11201\ : Span4Mux_v
    port map (
            O => \N__49410\,
            I => \N__49407\
        );

    \I__11200\ : Odrv4
    port map (
            O => \N__49407\,
            I => \pwm_generator_inst.un14_counter_5\
        );

    \I__11199\ : InMux
    port map (
            O => \N__49404\,
            I => \pwm_generator_inst.un19_threshold_0_cry_4\
        );

    \I__11198\ : CascadeMux
    port map (
            O => \N__49401\,
            I => \N__49398\
        );

    \I__11197\ : InMux
    port map (
            O => \N__49398\,
            I => \N__49395\
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__49395\,
            I => \N__49392\
        );

    \I__11195\ : Span4Mux_h
    port map (
            O => \N__49392\,
            I => \N__49389\
        );

    \I__11194\ : Odrv4
    port map (
            O => \N__49389\,
            I => \pwm_generator_inst.un14_counter_6\
        );

    \I__11193\ : InMux
    port map (
            O => \N__49386\,
            I => \pwm_generator_inst.un19_threshold_0_cry_5\
        );

    \I__11192\ : InMux
    port map (
            O => \N__49383\,
            I => \N__49379\
        );

    \I__11191\ : InMux
    port map (
            O => \N__49382\,
            I => \N__49375\
        );

    \I__11190\ : LocalMux
    port map (
            O => \N__49379\,
            I => \N__49372\
        );

    \I__11189\ : InMux
    port map (
            O => \N__49378\,
            I => \N__49369\
        );

    \I__11188\ : LocalMux
    port map (
            O => \N__49375\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__11187\ : Odrv4
    port map (
            O => \N__49372\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__11186\ : LocalMux
    port map (
            O => \N__49369\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__11185\ : InMux
    port map (
            O => \N__49362\,
            I => \N__49359\
        );

    \I__11184\ : LocalMux
    port map (
            O => \N__49359\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__11183\ : InMux
    port map (
            O => \N__49356\,
            I => \N__49352\
        );

    \I__11182\ : InMux
    port map (
            O => \N__49355\,
            I => \N__49348\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__49352\,
            I => \N__49345\
        );

    \I__11180\ : InMux
    port map (
            O => \N__49351\,
            I => \N__49342\
        );

    \I__11179\ : LocalMux
    port map (
            O => \N__49348\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__11178\ : Odrv4
    port map (
            O => \N__49345\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__11177\ : LocalMux
    port map (
            O => \N__49342\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__11176\ : InMux
    port map (
            O => \N__49335\,
            I => \N__49332\
        );

    \I__11175\ : LocalMux
    port map (
            O => \N__49332\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__11174\ : InMux
    port map (
            O => \N__49329\,
            I => \N__49325\
        );

    \I__11173\ : InMux
    port map (
            O => \N__49328\,
            I => \N__49321\
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__49325\,
            I => \N__49318\
        );

    \I__11171\ : InMux
    port map (
            O => \N__49324\,
            I => \N__49315\
        );

    \I__11170\ : LocalMux
    port map (
            O => \N__49321\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__11169\ : Odrv4
    port map (
            O => \N__49318\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__49315\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__11167\ : InMux
    port map (
            O => \N__49308\,
            I => \N__49305\
        );

    \I__11166\ : LocalMux
    port map (
            O => \N__49305\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__11165\ : InMux
    port map (
            O => \N__49302\,
            I => \N__49298\
        );

    \I__11164\ : InMux
    port map (
            O => \N__49301\,
            I => \N__49294\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__49298\,
            I => \N__49291\
        );

    \I__11162\ : InMux
    port map (
            O => \N__49297\,
            I => \N__49288\
        );

    \I__11161\ : LocalMux
    port map (
            O => \N__49294\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__11160\ : Odrv4
    port map (
            O => \N__49291\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__49288\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__11158\ : InMux
    port map (
            O => \N__49281\,
            I => \N__49278\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__49278\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__11156\ : InMux
    port map (
            O => \N__49275\,
            I => \N__49272\
        );

    \I__11155\ : LocalMux
    port map (
            O => \N__49272\,
            I => \N__49267\
        );

    \I__11154\ : InMux
    port map (
            O => \N__49271\,
            I => \N__49264\
        );

    \I__11153\ : InMux
    port map (
            O => \N__49270\,
            I => \N__49261\
        );

    \I__11152\ : Odrv4
    port map (
            O => \N__49267\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__11151\ : LocalMux
    port map (
            O => \N__49264\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__11150\ : LocalMux
    port map (
            O => \N__49261\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__11149\ : InMux
    port map (
            O => \N__49254\,
            I => \N__49251\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__49251\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__11147\ : InMux
    port map (
            O => \N__49248\,
            I => \N__49244\
        );

    \I__11146\ : InMux
    port map (
            O => \N__49247\,
            I => \N__49240\
        );

    \I__11145\ : LocalMux
    port map (
            O => \N__49244\,
            I => \N__49237\
        );

    \I__11144\ : InMux
    port map (
            O => \N__49243\,
            I => \N__49234\
        );

    \I__11143\ : LocalMux
    port map (
            O => \N__49240\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__11142\ : Odrv4
    port map (
            O => \N__49237\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__11141\ : LocalMux
    port map (
            O => \N__49234\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__11140\ : InMux
    port map (
            O => \N__49227\,
            I => \N__49224\
        );

    \I__11139\ : LocalMux
    port map (
            O => \N__49224\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__11138\ : InMux
    port map (
            O => \N__49221\,
            I => \N__49216\
        );

    \I__11137\ : InMux
    port map (
            O => \N__49220\,
            I => \N__49213\
        );

    \I__11136\ : InMux
    port map (
            O => \N__49219\,
            I => \N__49210\
        );

    \I__11135\ : LocalMux
    port map (
            O => \N__49216\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__11134\ : LocalMux
    port map (
            O => \N__49213\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__11133\ : LocalMux
    port map (
            O => \N__49210\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__11132\ : InMux
    port map (
            O => \N__49203\,
            I => \N__49200\
        );

    \I__11131\ : LocalMux
    port map (
            O => \N__49200\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__11130\ : InMux
    port map (
            O => \N__49197\,
            I => \N__49192\
        );

    \I__11129\ : InMux
    port map (
            O => \N__49196\,
            I => \N__49189\
        );

    \I__11128\ : InMux
    port map (
            O => \N__49195\,
            I => \N__49186\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__49192\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__49189\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__11125\ : LocalMux
    port map (
            O => \N__49186\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__11124\ : InMux
    port map (
            O => \N__49179\,
            I => \N__49176\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__49176\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__11122\ : CascadeMux
    port map (
            O => \N__49173\,
            I => \N__49170\
        );

    \I__11121\ : InMux
    port map (
            O => \N__49170\,
            I => \N__49167\
        );

    \I__11120\ : LocalMux
    port map (
            O => \N__49167\,
            I => \N__49162\
        );

    \I__11119\ : InMux
    port map (
            O => \N__49166\,
            I => \N__49159\
        );

    \I__11118\ : InMux
    port map (
            O => \N__49165\,
            I => \N__49156\
        );

    \I__11117\ : Span4Mux_h
    port map (
            O => \N__49162\,
            I => \N__49153\
        );

    \I__11116\ : LocalMux
    port map (
            O => \N__49159\,
            I => \N__49150\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__49156\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__11114\ : Odrv4
    port map (
            O => \N__49153\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__11113\ : Odrv12
    port map (
            O => \N__49150\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__11112\ : InMux
    port map (
            O => \N__49143\,
            I => \bfn_17_23_0_\
        );

    \I__11111\ : CascadeMux
    port map (
            O => \N__49140\,
            I => \N__49137\
        );

    \I__11110\ : InMux
    port map (
            O => \N__49137\,
            I => \N__49133\
        );

    \I__11109\ : CascadeMux
    port map (
            O => \N__49136\,
            I => \N__49130\
        );

    \I__11108\ : LocalMux
    port map (
            O => \N__49133\,
            I => \N__49126\
        );

    \I__11107\ : InMux
    port map (
            O => \N__49130\,
            I => \N__49123\
        );

    \I__11106\ : InMux
    port map (
            O => \N__49129\,
            I => \N__49120\
        );

    \I__11105\ : Span4Mux_h
    port map (
            O => \N__49126\,
            I => \N__49117\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__49123\,
            I => \N__49114\
        );

    \I__11103\ : LocalMux
    port map (
            O => \N__49120\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__11102\ : Odrv4
    port map (
            O => \N__49117\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__11101\ : Odrv12
    port map (
            O => \N__49114\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__11100\ : InMux
    port map (
            O => \N__49107\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__11099\ : InMux
    port map (
            O => \N__49104\,
            I => \N__49097\
        );

    \I__11098\ : InMux
    port map (
            O => \N__49103\,
            I => \N__49097\
        );

    \I__11097\ : InMux
    port map (
            O => \N__49102\,
            I => \N__49094\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__49097\,
            I => \N__49091\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__49094\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__11094\ : Odrv12
    port map (
            O => \N__49091\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__11093\ : InMux
    port map (
            O => \N__49086\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__11092\ : InMux
    port map (
            O => \N__49083\,
            I => \N__49076\
        );

    \I__11091\ : InMux
    port map (
            O => \N__49082\,
            I => \N__49076\
        );

    \I__11090\ : InMux
    port map (
            O => \N__49081\,
            I => \N__49073\
        );

    \I__11089\ : LocalMux
    port map (
            O => \N__49076\,
            I => \N__49070\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__49073\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__11087\ : Odrv12
    port map (
            O => \N__49070\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__11086\ : InMux
    port map (
            O => \N__49065\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__11085\ : CascadeMux
    port map (
            O => \N__49062\,
            I => \N__49059\
        );

    \I__11084\ : InMux
    port map (
            O => \N__49059\,
            I => \N__49055\
        );

    \I__11083\ : InMux
    port map (
            O => \N__49058\,
            I => \N__49052\
        );

    \I__11082\ : LocalMux
    port map (
            O => \N__49055\,
            I => \N__49049\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__49052\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__11080\ : Odrv12
    port map (
            O => \N__49049\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__11079\ : InMux
    port map (
            O => \N__49044\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__11078\ : InMux
    port map (
            O => \N__49041\,
            I => \N__49003\
        );

    \I__11077\ : InMux
    port map (
            O => \N__49040\,
            I => \N__49003\
        );

    \I__11076\ : InMux
    port map (
            O => \N__49039\,
            I => \N__49003\
        );

    \I__11075\ : InMux
    port map (
            O => \N__49038\,
            I => \N__49003\
        );

    \I__11074\ : InMux
    port map (
            O => \N__49037\,
            I => \N__48994\
        );

    \I__11073\ : InMux
    port map (
            O => \N__49036\,
            I => \N__48994\
        );

    \I__11072\ : InMux
    port map (
            O => \N__49035\,
            I => \N__48994\
        );

    \I__11071\ : InMux
    port map (
            O => \N__49034\,
            I => \N__48994\
        );

    \I__11070\ : InMux
    port map (
            O => \N__49033\,
            I => \N__48985\
        );

    \I__11069\ : InMux
    port map (
            O => \N__49032\,
            I => \N__48985\
        );

    \I__11068\ : InMux
    port map (
            O => \N__49031\,
            I => \N__48985\
        );

    \I__11067\ : InMux
    port map (
            O => \N__49030\,
            I => \N__48985\
        );

    \I__11066\ : InMux
    port map (
            O => \N__49029\,
            I => \N__48976\
        );

    \I__11065\ : InMux
    port map (
            O => \N__49028\,
            I => \N__48976\
        );

    \I__11064\ : InMux
    port map (
            O => \N__49027\,
            I => \N__48976\
        );

    \I__11063\ : InMux
    port map (
            O => \N__49026\,
            I => \N__48976\
        );

    \I__11062\ : InMux
    port map (
            O => \N__49025\,
            I => \N__48971\
        );

    \I__11061\ : InMux
    port map (
            O => \N__49024\,
            I => \N__48971\
        );

    \I__11060\ : InMux
    port map (
            O => \N__49023\,
            I => \N__48962\
        );

    \I__11059\ : InMux
    port map (
            O => \N__49022\,
            I => \N__48962\
        );

    \I__11058\ : InMux
    port map (
            O => \N__49021\,
            I => \N__48962\
        );

    \I__11057\ : InMux
    port map (
            O => \N__49020\,
            I => \N__48962\
        );

    \I__11056\ : InMux
    port map (
            O => \N__49019\,
            I => \N__48953\
        );

    \I__11055\ : InMux
    port map (
            O => \N__49018\,
            I => \N__48953\
        );

    \I__11054\ : InMux
    port map (
            O => \N__49017\,
            I => \N__48953\
        );

    \I__11053\ : InMux
    port map (
            O => \N__49016\,
            I => \N__48953\
        );

    \I__11052\ : InMux
    port map (
            O => \N__49015\,
            I => \N__48944\
        );

    \I__11051\ : InMux
    port map (
            O => \N__49014\,
            I => \N__48944\
        );

    \I__11050\ : InMux
    port map (
            O => \N__49013\,
            I => \N__48944\
        );

    \I__11049\ : InMux
    port map (
            O => \N__49012\,
            I => \N__48944\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__49003\,
            I => \N__48937\
        );

    \I__11047\ : LocalMux
    port map (
            O => \N__48994\,
            I => \N__48937\
        );

    \I__11046\ : LocalMux
    port map (
            O => \N__48985\,
            I => \N__48937\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__48976\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__11044\ : LocalMux
    port map (
            O => \N__48971\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__48962\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__11042\ : LocalMux
    port map (
            O => \N__48953\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__11041\ : LocalMux
    port map (
            O => \N__48944\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__11040\ : Odrv4
    port map (
            O => \N__48937\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__11039\ : InMux
    port map (
            O => \N__48924\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__11038\ : CascadeMux
    port map (
            O => \N__48921\,
            I => \N__48918\
        );

    \I__11037\ : InMux
    port map (
            O => \N__48918\,
            I => \N__48914\
        );

    \I__11036\ : InMux
    port map (
            O => \N__48917\,
            I => \N__48911\
        );

    \I__11035\ : LocalMux
    port map (
            O => \N__48914\,
            I => \N__48908\
        );

    \I__11034\ : LocalMux
    port map (
            O => \N__48911\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__11033\ : Odrv12
    port map (
            O => \N__48908\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__11032\ : CEMux
    port map (
            O => \N__48903\,
            I => \N__48899\
        );

    \I__11031\ : CEMux
    port map (
            O => \N__48902\,
            I => \N__48895\
        );

    \I__11030\ : LocalMux
    port map (
            O => \N__48899\,
            I => \N__48892\
        );

    \I__11029\ : CEMux
    port map (
            O => \N__48898\,
            I => \N__48889\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__48895\,
            I => \N__48885\
        );

    \I__11027\ : Span4Mux_v
    port map (
            O => \N__48892\,
            I => \N__48882\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__48889\,
            I => \N__48879\
        );

    \I__11025\ : CEMux
    port map (
            O => \N__48888\,
            I => \N__48876\
        );

    \I__11024\ : Span4Mux_h
    port map (
            O => \N__48885\,
            I => \N__48873\
        );

    \I__11023\ : Span4Mux_h
    port map (
            O => \N__48882\,
            I => \N__48870\
        );

    \I__11022\ : Span4Mux_h
    port map (
            O => \N__48879\,
            I => \N__48867\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__48876\,
            I => \N__48864\
        );

    \I__11020\ : Odrv4
    port map (
            O => \N__48873\,
            I => \delay_measurement_inst.delay_hc_timer.N_156_i\
        );

    \I__11019\ : Odrv4
    port map (
            O => \N__48870\,
            I => \delay_measurement_inst.delay_hc_timer.N_156_i\
        );

    \I__11018\ : Odrv4
    port map (
            O => \N__48867\,
            I => \delay_measurement_inst.delay_hc_timer.N_156_i\
        );

    \I__11017\ : Odrv12
    port map (
            O => \N__48864\,
            I => \delay_measurement_inst.delay_hc_timer.N_156_i\
        );

    \I__11016\ : InMux
    port map (
            O => \N__48855\,
            I => \N__48850\
        );

    \I__11015\ : InMux
    port map (
            O => \N__48854\,
            I => \N__48847\
        );

    \I__11014\ : InMux
    port map (
            O => \N__48853\,
            I => \N__48844\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__48850\,
            I => \N__48841\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__48847\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__48844\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__11010\ : Odrv4
    port map (
            O => \N__48841\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__11009\ : InMux
    port map (
            O => \N__48834\,
            I => \N__48831\
        );

    \I__11008\ : LocalMux
    port map (
            O => \N__48831\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__11007\ : InMux
    port map (
            O => \N__48828\,
            I => \N__48823\
        );

    \I__11006\ : InMux
    port map (
            O => \N__48827\,
            I => \N__48820\
        );

    \I__11005\ : InMux
    port map (
            O => \N__48826\,
            I => \N__48817\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__48823\,
            I => \N__48814\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__48820\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__48817\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__11001\ : Odrv4
    port map (
            O => \N__48814\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__11000\ : InMux
    port map (
            O => \N__48807\,
            I => \N__48804\
        );

    \I__10999\ : LocalMux
    port map (
            O => \N__48804\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__10998\ : InMux
    port map (
            O => \N__48801\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__10997\ : CascadeMux
    port map (
            O => \N__48798\,
            I => \N__48794\
        );

    \I__10996\ : CascadeMux
    port map (
            O => \N__48797\,
            I => \N__48791\
        );

    \I__10995\ : InMux
    port map (
            O => \N__48794\,
            I => \N__48788\
        );

    \I__10994\ : InMux
    port map (
            O => \N__48791\,
            I => \N__48785\
        );

    \I__10993\ : LocalMux
    port map (
            O => \N__48788\,
            I => \N__48779\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__48785\,
            I => \N__48779\
        );

    \I__10991\ : InMux
    port map (
            O => \N__48784\,
            I => \N__48776\
        );

    \I__10990\ : Span4Mux_v
    port map (
            O => \N__48779\,
            I => \N__48773\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__48776\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__10988\ : Odrv4
    port map (
            O => \N__48773\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__10987\ : InMux
    port map (
            O => \N__48768\,
            I => \bfn_17_22_0_\
        );

    \I__10986\ : CascadeMux
    port map (
            O => \N__48765\,
            I => \N__48761\
        );

    \I__10985\ : InMux
    port map (
            O => \N__48764\,
            I => \N__48758\
        );

    \I__10984\ : InMux
    port map (
            O => \N__48761\,
            I => \N__48755\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__48758\,
            I => \N__48751\
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__48755\,
            I => \N__48748\
        );

    \I__10981\ : InMux
    port map (
            O => \N__48754\,
            I => \N__48745\
        );

    \I__10980\ : Span4Mux_v
    port map (
            O => \N__48751\,
            I => \N__48740\
        );

    \I__10979\ : Span4Mux_v
    port map (
            O => \N__48748\,
            I => \N__48740\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__48745\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__10977\ : Odrv4
    port map (
            O => \N__48740\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__10976\ : InMux
    port map (
            O => \N__48735\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__10975\ : CascadeMux
    port map (
            O => \N__48732\,
            I => \N__48729\
        );

    \I__10974\ : InMux
    port map (
            O => \N__48729\,
            I => \N__48725\
        );

    \I__10973\ : InMux
    port map (
            O => \N__48728\,
            I => \N__48722\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__48725\,
            I => \N__48716\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__48722\,
            I => \N__48716\
        );

    \I__10970\ : InMux
    port map (
            O => \N__48721\,
            I => \N__48713\
        );

    \I__10969\ : Span4Mux_h
    port map (
            O => \N__48716\,
            I => \N__48710\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__48713\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__10967\ : Odrv4
    port map (
            O => \N__48710\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__10966\ : InMux
    port map (
            O => \N__48705\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__10965\ : CascadeMux
    port map (
            O => \N__48702\,
            I => \N__48698\
        );

    \I__10964\ : CascadeMux
    port map (
            O => \N__48701\,
            I => \N__48695\
        );

    \I__10963\ : InMux
    port map (
            O => \N__48698\,
            I => \N__48689\
        );

    \I__10962\ : InMux
    port map (
            O => \N__48695\,
            I => \N__48689\
        );

    \I__10961\ : InMux
    port map (
            O => \N__48694\,
            I => \N__48686\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__48689\,
            I => \N__48683\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__48686\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__10958\ : Odrv12
    port map (
            O => \N__48683\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__10957\ : InMux
    port map (
            O => \N__48678\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__10956\ : InMux
    port map (
            O => \N__48675\,
            I => \N__48668\
        );

    \I__10955\ : InMux
    port map (
            O => \N__48674\,
            I => \N__48668\
        );

    \I__10954\ : InMux
    port map (
            O => \N__48673\,
            I => \N__48665\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__48668\,
            I => \N__48662\
        );

    \I__10952\ : LocalMux
    port map (
            O => \N__48665\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__10951\ : Odrv12
    port map (
            O => \N__48662\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__10950\ : InMux
    port map (
            O => \N__48657\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__10949\ : CascadeMux
    port map (
            O => \N__48654\,
            I => \N__48651\
        );

    \I__10948\ : InMux
    port map (
            O => \N__48651\,
            I => \N__48646\
        );

    \I__10947\ : InMux
    port map (
            O => \N__48650\,
            I => \N__48643\
        );

    \I__10946\ : InMux
    port map (
            O => \N__48649\,
            I => \N__48640\
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__48646\,
            I => \N__48635\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__48643\,
            I => \N__48635\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__48640\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__10942\ : Odrv12
    port map (
            O => \N__48635\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__10941\ : InMux
    port map (
            O => \N__48630\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__10940\ : CascadeMux
    port map (
            O => \N__48627\,
            I => \N__48623\
        );

    \I__10939\ : CascadeMux
    port map (
            O => \N__48626\,
            I => \N__48620\
        );

    \I__10938\ : InMux
    port map (
            O => \N__48623\,
            I => \N__48614\
        );

    \I__10937\ : InMux
    port map (
            O => \N__48620\,
            I => \N__48614\
        );

    \I__10936\ : InMux
    port map (
            O => \N__48619\,
            I => \N__48611\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__48614\,
            I => \N__48608\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__48611\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__10933\ : Odrv12
    port map (
            O => \N__48608\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__10932\ : InMux
    port map (
            O => \N__48603\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__10931\ : InMux
    port map (
            O => \N__48600\,
            I => \N__48593\
        );

    \I__10930\ : InMux
    port map (
            O => \N__48599\,
            I => \N__48593\
        );

    \I__10929\ : InMux
    port map (
            O => \N__48598\,
            I => \N__48590\
        );

    \I__10928\ : LocalMux
    port map (
            O => \N__48593\,
            I => \N__48587\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__48590\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__10926\ : Odrv12
    port map (
            O => \N__48587\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__10925\ : InMux
    port map (
            O => \N__48582\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__10924\ : CascadeMux
    port map (
            O => \N__48579\,
            I => \N__48575\
        );

    \I__10923\ : CascadeMux
    port map (
            O => \N__48578\,
            I => \N__48572\
        );

    \I__10922\ : InMux
    port map (
            O => \N__48575\,
            I => \N__48567\
        );

    \I__10921\ : InMux
    port map (
            O => \N__48572\,
            I => \N__48567\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__48567\,
            I => \N__48563\
        );

    \I__10919\ : InMux
    port map (
            O => \N__48566\,
            I => \N__48560\
        );

    \I__10918\ : Span4Mux_v
    port map (
            O => \N__48563\,
            I => \N__48557\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__48560\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__10916\ : Odrv4
    port map (
            O => \N__48557\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__10915\ : InMux
    port map (
            O => \N__48552\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__10914\ : CascadeMux
    port map (
            O => \N__48549\,
            I => \N__48546\
        );

    \I__10913\ : InMux
    port map (
            O => \N__48546\,
            I => \N__48543\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__48543\,
            I => \N__48538\
        );

    \I__10911\ : InMux
    port map (
            O => \N__48542\,
            I => \N__48535\
        );

    \I__10910\ : InMux
    port map (
            O => \N__48541\,
            I => \N__48532\
        );

    \I__10909\ : Span4Mux_h
    port map (
            O => \N__48538\,
            I => \N__48529\
        );

    \I__10908\ : LocalMux
    port map (
            O => \N__48535\,
            I => \N__48526\
        );

    \I__10907\ : LocalMux
    port map (
            O => \N__48532\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__10906\ : Odrv4
    port map (
            O => \N__48529\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__10905\ : Odrv12
    port map (
            O => \N__48526\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__10904\ : InMux
    port map (
            O => \N__48519\,
            I => \bfn_17_21_0_\
        );

    \I__10903\ : CascadeMux
    port map (
            O => \N__48516\,
            I => \N__48513\
        );

    \I__10902\ : InMux
    port map (
            O => \N__48513\,
            I => \N__48509\
        );

    \I__10901\ : InMux
    port map (
            O => \N__48512\,
            I => \N__48506\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__48509\,
            I => \N__48500\
        );

    \I__10899\ : LocalMux
    port map (
            O => \N__48506\,
            I => \N__48500\
        );

    \I__10898\ : InMux
    port map (
            O => \N__48505\,
            I => \N__48497\
        );

    \I__10897\ : Span4Mux_v
    port map (
            O => \N__48500\,
            I => \N__48494\
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__48497\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__10895\ : Odrv4
    port map (
            O => \N__48494\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__10894\ : InMux
    port map (
            O => \N__48489\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__10893\ : InMux
    port map (
            O => \N__48486\,
            I => \N__48480\
        );

    \I__10892\ : InMux
    port map (
            O => \N__48485\,
            I => \N__48480\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__48480\,
            I => \N__48476\
        );

    \I__10890\ : InMux
    port map (
            O => \N__48479\,
            I => \N__48473\
        );

    \I__10889\ : Span4Mux_h
    port map (
            O => \N__48476\,
            I => \N__48470\
        );

    \I__10888\ : LocalMux
    port map (
            O => \N__48473\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__10887\ : Odrv4
    port map (
            O => \N__48470\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__10886\ : InMux
    port map (
            O => \N__48465\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__10885\ : InMux
    port map (
            O => \N__48462\,
            I => \N__48456\
        );

    \I__10884\ : InMux
    port map (
            O => \N__48461\,
            I => \N__48456\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__48456\,
            I => \N__48452\
        );

    \I__10882\ : InMux
    port map (
            O => \N__48455\,
            I => \N__48449\
        );

    \I__10881\ : Span4Mux_h
    port map (
            O => \N__48452\,
            I => \N__48446\
        );

    \I__10880\ : LocalMux
    port map (
            O => \N__48449\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__10879\ : Odrv4
    port map (
            O => \N__48446\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__10878\ : InMux
    port map (
            O => \N__48441\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__10877\ : CascadeMux
    port map (
            O => \N__48438\,
            I => \N__48434\
        );

    \I__10876\ : CascadeMux
    port map (
            O => \N__48437\,
            I => \N__48431\
        );

    \I__10875\ : InMux
    port map (
            O => \N__48434\,
            I => \N__48426\
        );

    \I__10874\ : InMux
    port map (
            O => \N__48431\,
            I => \N__48426\
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__48426\,
            I => \N__48422\
        );

    \I__10872\ : InMux
    port map (
            O => \N__48425\,
            I => \N__48419\
        );

    \I__10871\ : Span4Mux_v
    port map (
            O => \N__48422\,
            I => \N__48416\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__48419\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__10869\ : Odrv4
    port map (
            O => \N__48416\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__10868\ : InMux
    port map (
            O => \N__48411\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__10867\ : CascadeMux
    port map (
            O => \N__48408\,
            I => \N__48404\
        );

    \I__10866\ : CascadeMux
    port map (
            O => \N__48407\,
            I => \N__48401\
        );

    \I__10865\ : InMux
    port map (
            O => \N__48404\,
            I => \N__48396\
        );

    \I__10864\ : InMux
    port map (
            O => \N__48401\,
            I => \N__48396\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__48396\,
            I => \N__48392\
        );

    \I__10862\ : InMux
    port map (
            O => \N__48395\,
            I => \N__48389\
        );

    \I__10861\ : Span4Mux_h
    port map (
            O => \N__48392\,
            I => \N__48386\
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__48389\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__10859\ : Odrv4
    port map (
            O => \N__48386\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__10858\ : InMux
    port map (
            O => \N__48381\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__10857\ : InMux
    port map (
            O => \N__48378\,
            I => \N__48372\
        );

    \I__10856\ : InMux
    port map (
            O => \N__48377\,
            I => \N__48372\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__48372\,
            I => \N__48368\
        );

    \I__10854\ : InMux
    port map (
            O => \N__48371\,
            I => \N__48365\
        );

    \I__10853\ : Span4Mux_v
    port map (
            O => \N__48368\,
            I => \N__48362\
        );

    \I__10852\ : LocalMux
    port map (
            O => \N__48365\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__10851\ : Odrv4
    port map (
            O => \N__48362\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__10850\ : InMux
    port map (
            O => \N__48357\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__10849\ : InMux
    port map (
            O => \N__48354\,
            I => \N__48348\
        );

    \I__10848\ : InMux
    port map (
            O => \N__48353\,
            I => \N__48348\
        );

    \I__10847\ : LocalMux
    port map (
            O => \N__48348\,
            I => \N__48344\
        );

    \I__10846\ : InMux
    port map (
            O => \N__48347\,
            I => \N__48341\
        );

    \I__10845\ : Span4Mux_v
    port map (
            O => \N__48344\,
            I => \N__48338\
        );

    \I__10844\ : LocalMux
    port map (
            O => \N__48341\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__10843\ : Odrv4
    port map (
            O => \N__48338\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__10842\ : InMux
    port map (
            O => \N__48333\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__10841\ : InMux
    port map (
            O => \N__48330\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__10840\ : InMux
    port map (
            O => \N__48327\,
            I => \N__48323\
        );

    \I__10839\ : InMux
    port map (
            O => \N__48326\,
            I => \N__48320\
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__48323\,
            I => \N__48317\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__48320\,
            I => \N__48314\
        );

    \I__10836\ : Span4Mux_h
    port map (
            O => \N__48317\,
            I => \N__48309\
        );

    \I__10835\ : Span4Mux_h
    port map (
            O => \N__48314\,
            I => \N__48309\
        );

    \I__10834\ : Odrv4
    port map (
            O => \N__48309\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__10833\ : InMux
    port map (
            O => \N__48306\,
            I => \bfn_17_20_0_\
        );

    \I__10832\ : InMux
    port map (
            O => \N__48303\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__10831\ : InMux
    port map (
            O => \N__48300\,
            I => \N__48293\
        );

    \I__10830\ : InMux
    port map (
            O => \N__48299\,
            I => \N__48293\
        );

    \I__10829\ : InMux
    port map (
            O => \N__48298\,
            I => \N__48290\
        );

    \I__10828\ : LocalMux
    port map (
            O => \N__48293\,
            I => \N__48287\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__48290\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__10826\ : Odrv12
    port map (
            O => \N__48287\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__10825\ : InMux
    port map (
            O => \N__48282\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__10824\ : InMux
    port map (
            O => \N__48279\,
            I => \N__48272\
        );

    \I__10823\ : InMux
    port map (
            O => \N__48278\,
            I => \N__48272\
        );

    \I__10822\ : InMux
    port map (
            O => \N__48277\,
            I => \N__48269\
        );

    \I__10821\ : LocalMux
    port map (
            O => \N__48272\,
            I => \N__48266\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__48269\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__10819\ : Odrv12
    port map (
            O => \N__48266\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__10818\ : InMux
    port map (
            O => \N__48261\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__10817\ : CascadeMux
    port map (
            O => \N__48258\,
            I => \N__48254\
        );

    \I__10816\ : InMux
    port map (
            O => \N__48257\,
            I => \N__48250\
        );

    \I__10815\ : InMux
    port map (
            O => \N__48254\,
            I => \N__48247\
        );

    \I__10814\ : InMux
    port map (
            O => \N__48253\,
            I => \N__48244\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__48250\,
            I => \N__48239\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__48247\,
            I => \N__48239\
        );

    \I__10811\ : LocalMux
    port map (
            O => \N__48244\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__10810\ : Odrv12
    port map (
            O => \N__48239\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__10809\ : InMux
    port map (
            O => \N__48234\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__10808\ : CascadeMux
    port map (
            O => \N__48231\,
            I => \N__48227\
        );

    \I__10807\ : InMux
    port map (
            O => \N__48230\,
            I => \N__48224\
        );

    \I__10806\ : InMux
    port map (
            O => \N__48227\,
            I => \N__48221\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__48224\,
            I => \N__48217\
        );

    \I__10804\ : LocalMux
    port map (
            O => \N__48221\,
            I => \N__48214\
        );

    \I__10803\ : InMux
    port map (
            O => \N__48220\,
            I => \N__48211\
        );

    \I__10802\ : Span4Mux_h
    port map (
            O => \N__48217\,
            I => \N__48206\
        );

    \I__10801\ : Span4Mux_h
    port map (
            O => \N__48214\,
            I => \N__48206\
        );

    \I__10800\ : LocalMux
    port map (
            O => \N__48211\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__10799\ : Odrv4
    port map (
            O => \N__48206\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__10798\ : InMux
    port map (
            O => \N__48201\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__10797\ : CascadeMux
    port map (
            O => \N__48198\,
            I => \N__48194\
        );

    \I__10796\ : CascadeMux
    port map (
            O => \N__48197\,
            I => \N__48191\
        );

    \I__10795\ : InMux
    port map (
            O => \N__48194\,
            I => \N__48186\
        );

    \I__10794\ : InMux
    port map (
            O => \N__48191\,
            I => \N__48186\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__48186\,
            I => \N__48182\
        );

    \I__10792\ : InMux
    port map (
            O => \N__48185\,
            I => \N__48179\
        );

    \I__10791\ : Span4Mux_v
    port map (
            O => \N__48182\,
            I => \N__48176\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__48179\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__10789\ : Odrv4
    port map (
            O => \N__48176\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__10788\ : InMux
    port map (
            O => \N__48171\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__10787\ : InMux
    port map (
            O => \N__48168\,
            I => \N__48164\
        );

    \I__10786\ : CascadeMux
    port map (
            O => \N__48167\,
            I => \N__48161\
        );

    \I__10785\ : LocalMux
    port map (
            O => \N__48164\,
            I => \N__48158\
        );

    \I__10784\ : InMux
    port map (
            O => \N__48161\,
            I => \N__48155\
        );

    \I__10783\ : Odrv4
    port map (
            O => \N__48158\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__48155\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__10781\ : InMux
    port map (
            O => \N__48150\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__10780\ : InMux
    port map (
            O => \N__48147\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__10779\ : InMux
    port map (
            O => \N__48144\,
            I => \N__48141\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__48141\,
            I => \N__48138\
        );

    \I__10777\ : Span4Mux_h
    port map (
            O => \N__48138\,
            I => \N__48134\
        );

    \I__10776\ : InMux
    port map (
            O => \N__48137\,
            I => \N__48131\
        );

    \I__10775\ : Odrv4
    port map (
            O => \N__48134\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__48131\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__10773\ : InMux
    port map (
            O => \N__48126\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__10772\ : CascadeMux
    port map (
            O => \N__48123\,
            I => \N__48119\
        );

    \I__10771\ : InMux
    port map (
            O => \N__48122\,
            I => \N__48114\
        );

    \I__10770\ : InMux
    port map (
            O => \N__48119\,
            I => \N__48114\
        );

    \I__10769\ : LocalMux
    port map (
            O => \N__48114\,
            I => \N__48111\
        );

    \I__10768\ : Odrv4
    port map (
            O => \N__48111\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__10767\ : InMux
    port map (
            O => \N__48108\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__10766\ : InMux
    port map (
            O => \N__48105\,
            I => \N__48099\
        );

    \I__10765\ : InMux
    port map (
            O => \N__48104\,
            I => \N__48099\
        );

    \I__10764\ : LocalMux
    port map (
            O => \N__48099\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__10763\ : InMux
    port map (
            O => \N__48096\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__10762\ : InMux
    port map (
            O => \N__48093\,
            I => \bfn_17_19_0_\
        );

    \I__10761\ : InMux
    port map (
            O => \N__48090\,
            I => \N__48087\
        );

    \I__10760\ : LocalMux
    port map (
            O => \N__48087\,
            I => \N__48084\
        );

    \I__10759\ : Span4Mux_v
    port map (
            O => \N__48084\,
            I => \N__48081\
        );

    \I__10758\ : Span4Mux_v
    port map (
            O => \N__48081\,
            I => \N__48077\
        );

    \I__10757\ : InMux
    port map (
            O => \N__48080\,
            I => \N__48074\
        );

    \I__10756\ : Odrv4
    port map (
            O => \N__48077\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__10755\ : LocalMux
    port map (
            O => \N__48074\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__10754\ : InMux
    port map (
            O => \N__48069\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__10753\ : InMux
    port map (
            O => \N__48066\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__10752\ : InMux
    port map (
            O => \N__48063\,
            I => \N__48060\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__48060\,
            I => \N__48056\
        );

    \I__10750\ : CascadeMux
    port map (
            O => \N__48059\,
            I => \N__48053\
        );

    \I__10749\ : Span4Mux_h
    port map (
            O => \N__48056\,
            I => \N__48050\
        );

    \I__10748\ : InMux
    port map (
            O => \N__48053\,
            I => \N__48047\
        );

    \I__10747\ : Odrv4
    port map (
            O => \N__48050\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__10746\ : LocalMux
    port map (
            O => \N__48047\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__10745\ : InMux
    port map (
            O => \N__48042\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__10744\ : InMux
    port map (
            O => \N__48039\,
            I => \N__48036\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__48036\,
            I => \N__48033\
        );

    \I__10742\ : Span4Mux_h
    port map (
            O => \N__48033\,
            I => \N__48029\
        );

    \I__10741\ : InMux
    port map (
            O => \N__48032\,
            I => \N__48026\
        );

    \I__10740\ : Odrv4
    port map (
            O => \N__48029\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__48026\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__10738\ : InMux
    port map (
            O => \N__48021\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__10737\ : InMux
    port map (
            O => \N__48018\,
            I => \N__48015\
        );

    \I__10736\ : LocalMux
    port map (
            O => \N__48015\,
            I => \N__48011\
        );

    \I__10735\ : InMux
    port map (
            O => \N__48014\,
            I => \N__48008\
        );

    \I__10734\ : Odrv4
    port map (
            O => \N__48011\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__48008\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__10732\ : InMux
    port map (
            O => \N__48003\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__10731\ : InMux
    port map (
            O => \N__48000\,
            I => \N__47997\
        );

    \I__10730\ : LocalMux
    port map (
            O => \N__47997\,
            I => \N__47994\
        );

    \I__10729\ : Span4Mux_h
    port map (
            O => \N__47994\,
            I => \N__47990\
        );

    \I__10728\ : InMux
    port map (
            O => \N__47993\,
            I => \N__47987\
        );

    \I__10727\ : Odrv4
    port map (
            O => \N__47990\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__47987\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__10725\ : InMux
    port map (
            O => \N__47982\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__10724\ : InMux
    port map (
            O => \N__47979\,
            I => \N__47976\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__47976\,
            I => \N__47972\
        );

    \I__10722\ : InMux
    port map (
            O => \N__47975\,
            I => \N__47969\
        );

    \I__10721\ : Odrv4
    port map (
            O => \N__47972\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__47969\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10719\ : InMux
    port map (
            O => \N__47964\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__10718\ : InMux
    port map (
            O => \N__47961\,
            I => \N__47958\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__47958\,
            I => \N__47954\
        );

    \I__10716\ : CascadeMux
    port map (
            O => \N__47957\,
            I => \N__47951\
        );

    \I__10715\ : Span4Mux_v
    port map (
            O => \N__47954\,
            I => \N__47948\
        );

    \I__10714\ : InMux
    port map (
            O => \N__47951\,
            I => \N__47945\
        );

    \I__10713\ : Odrv4
    port map (
            O => \N__47948\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__47945\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__10711\ : InMux
    port map (
            O => \N__47940\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__10710\ : InMux
    port map (
            O => \N__47937\,
            I => \N__47934\
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__47934\,
            I => \N__47931\
        );

    \I__10708\ : Span4Mux_h
    port map (
            O => \N__47931\,
            I => \N__47927\
        );

    \I__10707\ : InMux
    port map (
            O => \N__47930\,
            I => \N__47924\
        );

    \I__10706\ : Odrv4
    port map (
            O => \N__47927\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__47924\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__10704\ : InMux
    port map (
            O => \N__47919\,
            I => \bfn_17_18_0_\
        );

    \I__10703\ : InMux
    port map (
            O => \N__47916\,
            I => \N__47913\
        );

    \I__10702\ : LocalMux
    port map (
            O => \N__47913\,
            I => \N__47910\
        );

    \I__10701\ : Span4Mux_h
    port map (
            O => \N__47910\,
            I => \N__47906\
        );

    \I__10700\ : InMux
    port map (
            O => \N__47909\,
            I => \N__47903\
        );

    \I__10699\ : Odrv4
    port map (
            O => \N__47906\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__10698\ : LocalMux
    port map (
            O => \N__47903\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__10697\ : InMux
    port map (
            O => \N__47898\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__10696\ : InMux
    port map (
            O => \N__47895\,
            I => \N__47891\
        );

    \I__10695\ : InMux
    port map (
            O => \N__47894\,
            I => \N__47888\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__47891\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__47888\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__10692\ : InMux
    port map (
            O => \N__47883\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__10691\ : InMux
    port map (
            O => \N__47880\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__10690\ : InMux
    port map (
            O => \N__47877\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__10689\ : InMux
    port map (
            O => \N__47874\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__10688\ : InMux
    port map (
            O => \N__47871\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__10687\ : InMux
    port map (
            O => \N__47868\,
            I => \N__47865\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__47865\,
            I => \N__47862\
        );

    \I__10685\ : Span4Mux_h
    port map (
            O => \N__47862\,
            I => \N__47858\
        );

    \I__10684\ : InMux
    port map (
            O => \N__47861\,
            I => \N__47855\
        );

    \I__10683\ : Odrv4
    port map (
            O => \N__47858\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__47855\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__10681\ : InMux
    port map (
            O => \N__47850\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__10680\ : InMux
    port map (
            O => \N__47847\,
            I => \N__47844\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__47844\,
            I => \N__47841\
        );

    \I__10678\ : Span4Mux_h
    port map (
            O => \N__47841\,
            I => \N__47837\
        );

    \I__10677\ : InMux
    port map (
            O => \N__47840\,
            I => \N__47834\
        );

    \I__10676\ : Odrv4
    port map (
            O => \N__47837\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__10675\ : LocalMux
    port map (
            O => \N__47834\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__10674\ : InMux
    port map (
            O => \N__47829\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__10673\ : InMux
    port map (
            O => \N__47826\,
            I => \N__47823\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__47823\,
            I => \N__47819\
        );

    \I__10671\ : InMux
    port map (
            O => \N__47822\,
            I => \N__47816\
        );

    \I__10670\ : Odrv4
    port map (
            O => \N__47819\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__10669\ : LocalMux
    port map (
            O => \N__47816\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__10668\ : InMux
    port map (
            O => \N__47811\,
            I => \bfn_17_17_0_\
        );

    \I__10667\ : InMux
    port map (
            O => \N__47808\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__10666\ : InMux
    port map (
            O => \N__47805\,
            I => \N__47802\
        );

    \I__10665\ : LocalMux
    port map (
            O => \N__47802\,
            I => \N__47799\
        );

    \I__10664\ : Odrv4
    port map (
            O => \N__47799\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26\
        );

    \I__10663\ : InMux
    port map (
            O => \N__47796\,
            I => \N__47792\
        );

    \I__10662\ : InMux
    port map (
            O => \N__47795\,
            I => \N__47789\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__47792\,
            I => \N__47784\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__47789\,
            I => \N__47784\
        );

    \I__10659\ : Span4Mux_v
    port map (
            O => \N__47784\,
            I => \N__47781\
        );

    \I__10658\ : Odrv4
    port map (
            O => \N__47781\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0\
        );

    \I__10657\ : InMux
    port map (
            O => \N__47778\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25\
        );

    \I__10656\ : InMux
    port map (
            O => \N__47775\,
            I => \N__47771\
        );

    \I__10655\ : InMux
    port map (
            O => \N__47774\,
            I => \N__47768\
        );

    \I__10654\ : LocalMux
    port map (
            O => \N__47771\,
            I => \N__47763\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__47768\,
            I => \N__47763\
        );

    \I__10652\ : Odrv12
    port map (
            O => \N__47763\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0\
        );

    \I__10651\ : InMux
    port map (
            O => \N__47760\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26\
        );

    \I__10650\ : InMux
    port map (
            O => \N__47757\,
            I => \N__47754\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__47754\,
            I => \N__47751\
        );

    \I__10648\ : Span4Mux_v
    port map (
            O => \N__47751\,
            I => \N__47748\
        );

    \I__10647\ : Odrv4
    port map (
            O => \N__47748\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28\
        );

    \I__10646\ : InMux
    port map (
            O => \N__47745\,
            I => \N__47741\
        );

    \I__10645\ : InMux
    port map (
            O => \N__47744\,
            I => \N__47738\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__47741\,
            I => \N__47733\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__47738\,
            I => \N__47733\
        );

    \I__10642\ : Odrv12
    port map (
            O => \N__47733\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0\
        );

    \I__10641\ : InMux
    port map (
            O => \N__47730\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27\
        );

    \I__10640\ : InMux
    port map (
            O => \N__47727\,
            I => \N__47723\
        );

    \I__10639\ : InMux
    port map (
            O => \N__47726\,
            I => \N__47720\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__47723\,
            I => \N__47715\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__47720\,
            I => \N__47715\
        );

    \I__10636\ : Span4Mux_v
    port map (
            O => \N__47715\,
            I => \N__47712\
        );

    \I__10635\ : Odrv4
    port map (
            O => \N__47712\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0\
        );

    \I__10634\ : InMux
    port map (
            O => \N__47709\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28\
        );

    \I__10633\ : InMux
    port map (
            O => \N__47706\,
            I => \N__47703\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__47703\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30\
        );

    \I__10631\ : InMux
    port map (
            O => \N__47700\,
            I => \N__47696\
        );

    \I__10630\ : InMux
    port map (
            O => \N__47699\,
            I => \N__47693\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__47696\,
            I => \N__47688\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__47693\,
            I => \N__47688\
        );

    \I__10627\ : Odrv12
    port map (
            O => \N__47688\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0\
        );

    \I__10626\ : InMux
    port map (
            O => \N__47685\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29\
        );

    \I__10625\ : InMux
    port map (
            O => \N__47682\,
            I => \N__47679\
        );

    \I__10624\ : LocalMux
    port map (
            O => \N__47679\,
            I => \N__47676\
        );

    \I__10623\ : Span4Mux_v
    port map (
            O => \N__47676\,
            I => \N__47673\
        );

    \I__10622\ : Odrv4
    port map (
            O => \N__47673\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO\
        );

    \I__10621\ : InMux
    port map (
            O => \N__47670\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30\
        );

    \I__10620\ : InMux
    port map (
            O => \N__47667\,
            I => \N__47664\
        );

    \I__10619\ : LocalMux
    port map (
            O => \N__47664\,
            I => \N__47661\
        );

    \I__10618\ : Span4Mux_h
    port map (
            O => \N__47661\,
            I => \N__47657\
        );

    \I__10617\ : InMux
    port map (
            O => \N__47660\,
            I => \N__47654\
        );

    \I__10616\ : Span4Mux_v
    port map (
            O => \N__47657\,
            I => \N__47651\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__47654\,
            I => \N__47648\
        );

    \I__10614\ : Odrv4
    port map (
            O => \N__47651\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_28
        );

    \I__10613\ : Odrv12
    port map (
            O => \N__47648\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_28
        );

    \I__10612\ : InMux
    port map (
            O => \N__47643\,
            I => \N__47639\
        );

    \I__10611\ : InMux
    port map (
            O => \N__47642\,
            I => \N__47636\
        );

    \I__10610\ : LocalMux
    port map (
            O => \N__47639\,
            I => \N__47632\
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__47636\,
            I => \N__47629\
        );

    \I__10608\ : InMux
    port map (
            O => \N__47635\,
            I => \N__47626\
        );

    \I__10607\ : Span4Mux_h
    port map (
            O => \N__47632\,
            I => \N__47622\
        );

    \I__10606\ : Span4Mux_h
    port map (
            O => \N__47629\,
            I => \N__47619\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__47626\,
            I => \N__47614\
        );

    \I__10604\ : InMux
    port map (
            O => \N__47625\,
            I => \N__47611\
        );

    \I__10603\ : Span4Mux_v
    port map (
            O => \N__47622\,
            I => \N__47608\
        );

    \I__10602\ : Span4Mux_h
    port map (
            O => \N__47619\,
            I => \N__47605\
        );

    \I__10601\ : InMux
    port map (
            O => \N__47618\,
            I => \N__47600\
        );

    \I__10600\ : InMux
    port map (
            O => \N__47617\,
            I => \N__47600\
        );

    \I__10599\ : Span12Mux_s9_v
    port map (
            O => \N__47614\,
            I => \N__47595\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__47611\,
            I => \N__47595\
        );

    \I__10597\ : Odrv4
    port map (
            O => \N__47608\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__10596\ : Odrv4
    port map (
            O => \N__47605\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__47600\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__10594\ : Odrv12
    port map (
            O => \N__47595\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__10593\ : InMux
    port map (
            O => \N__47586\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__10592\ : InMux
    port map (
            O => \N__47583\,
            I => \N__47580\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__47580\,
            I => \N__47577\
        );

    \I__10590\ : Odrv4
    port map (
            O => \N__47577\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18\
        );

    \I__10589\ : InMux
    port map (
            O => \N__47574\,
            I => \N__47570\
        );

    \I__10588\ : InMux
    port map (
            O => \N__47573\,
            I => \N__47567\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__47570\,
            I => \N__47562\
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__47567\,
            I => \N__47562\
        );

    \I__10585\ : Span4Mux_v
    port map (
            O => \N__47562\,
            I => \N__47559\
        );

    \I__10584\ : Odrv4
    port map (
            O => \N__47559\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9\
        );

    \I__10583\ : InMux
    port map (
            O => \N__47556\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17\
        );

    \I__10582\ : InMux
    port map (
            O => \N__47553\,
            I => \N__47550\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__47550\,
            I => \N__47547\
        );

    \I__10580\ : Span4Mux_h
    port map (
            O => \N__47547\,
            I => \N__47544\
        );

    \I__10579\ : Odrv4
    port map (
            O => \N__47544\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19\
        );

    \I__10578\ : InMux
    port map (
            O => \N__47541\,
            I => \N__47537\
        );

    \I__10577\ : InMux
    port map (
            O => \N__47540\,
            I => \N__47534\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__47537\,
            I => \N__47529\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__47534\,
            I => \N__47529\
        );

    \I__10574\ : Span4Mux_h
    port map (
            O => \N__47529\,
            I => \N__47526\
        );

    \I__10573\ : Odrv4
    port map (
            O => \N__47526\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9\
        );

    \I__10572\ : InMux
    port map (
            O => \N__47523\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18\
        );

    \I__10571\ : InMux
    port map (
            O => \N__47520\,
            I => \N__47517\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__47517\,
            I => \N__47514\
        );

    \I__10569\ : Odrv4
    port map (
            O => \N__47514\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20\
        );

    \I__10568\ : InMux
    port map (
            O => \N__47511\,
            I => \N__47507\
        );

    \I__10567\ : InMux
    port map (
            O => \N__47510\,
            I => \N__47504\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__47507\,
            I => \N__47499\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__47504\,
            I => \N__47499\
        );

    \I__10564\ : Span4Mux_h
    port map (
            O => \N__47499\,
            I => \N__47496\
        );

    \I__10563\ : Odrv4
    port map (
            O => \N__47496\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9\
        );

    \I__10562\ : InMux
    port map (
            O => \N__47493\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19\
        );

    \I__10561\ : InMux
    port map (
            O => \N__47490\,
            I => \N__47487\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__47487\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21\
        );

    \I__10559\ : InMux
    port map (
            O => \N__47484\,
            I => \N__47480\
        );

    \I__10558\ : InMux
    port map (
            O => \N__47483\,
            I => \N__47477\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__47480\,
            I => \N__47472\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__47477\,
            I => \N__47472\
        );

    \I__10555\ : Odrv12
    port map (
            O => \N__47472\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0\
        );

    \I__10554\ : InMux
    port map (
            O => \N__47469\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20\
        );

    \I__10553\ : InMux
    port map (
            O => \N__47466\,
            I => \N__47463\
        );

    \I__10552\ : LocalMux
    port map (
            O => \N__47463\,
            I => \N__47460\
        );

    \I__10551\ : Odrv4
    port map (
            O => \N__47460\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22\
        );

    \I__10550\ : InMux
    port map (
            O => \N__47457\,
            I => \N__47453\
        );

    \I__10549\ : InMux
    port map (
            O => \N__47456\,
            I => \N__47450\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__47453\,
            I => \N__47445\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__47450\,
            I => \N__47445\
        );

    \I__10546\ : Span4Mux_h
    port map (
            O => \N__47445\,
            I => \N__47442\
        );

    \I__10545\ : Odrv4
    port map (
            O => \N__47442\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0\
        );

    \I__10544\ : InMux
    port map (
            O => \N__47439\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21\
        );

    \I__10543\ : InMux
    port map (
            O => \N__47436\,
            I => \N__47432\
        );

    \I__10542\ : InMux
    port map (
            O => \N__47435\,
            I => \N__47429\
        );

    \I__10541\ : LocalMux
    port map (
            O => \N__47432\,
            I => \N__47424\
        );

    \I__10540\ : LocalMux
    port map (
            O => \N__47429\,
            I => \N__47424\
        );

    \I__10539\ : Odrv12
    port map (
            O => \N__47424\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0\
        );

    \I__10538\ : InMux
    port map (
            O => \N__47421\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22\
        );

    \I__10537\ : InMux
    port map (
            O => \N__47418\,
            I => \N__47415\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__47415\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24\
        );

    \I__10535\ : InMux
    port map (
            O => \N__47412\,
            I => \N__47408\
        );

    \I__10534\ : InMux
    port map (
            O => \N__47411\,
            I => \N__47405\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__47408\,
            I => \N__47400\
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__47405\,
            I => \N__47400\
        );

    \I__10531\ : Odrv12
    port map (
            O => \N__47400\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0\
        );

    \I__10530\ : InMux
    port map (
            O => \N__47397\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23\
        );

    \I__10529\ : InMux
    port map (
            O => \N__47394\,
            I => \N__47391\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__47391\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25\
        );

    \I__10527\ : InMux
    port map (
            O => \N__47388\,
            I => \N__47384\
        );

    \I__10526\ : InMux
    port map (
            O => \N__47387\,
            I => \N__47381\
        );

    \I__10525\ : LocalMux
    port map (
            O => \N__47384\,
            I => \N__47376\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__47381\,
            I => \N__47376\
        );

    \I__10523\ : Span4Mux_v
    port map (
            O => \N__47376\,
            I => \N__47373\
        );

    \I__10522\ : Odrv4
    port map (
            O => \N__47373\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0\
        );

    \I__10521\ : InMux
    port map (
            O => \N__47370\,
            I => \bfn_17_15_0_\
        );

    \I__10520\ : InMux
    port map (
            O => \N__47367\,
            I => \N__47364\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__47364\,
            I => \N__47360\
        );

    \I__10518\ : InMux
    port map (
            O => \N__47363\,
            I => \N__47357\
        );

    \I__10517\ : Span4Mux_v
    port map (
            O => \N__47360\,
            I => \N__47354\
        );

    \I__10516\ : LocalMux
    port map (
            O => \N__47357\,
            I => \N__47351\
        );

    \I__10515\ : Odrv4
    port map (
            O => \N__47354\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3\
        );

    \I__10514\ : Odrv12
    port map (
            O => \N__47351\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3\
        );

    \I__10513\ : InMux
    port map (
            O => \N__47346\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9\
        );

    \I__10512\ : InMux
    port map (
            O => \N__47343\,
            I => \N__47340\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__47340\,
            I => \N__47337\
        );

    \I__10510\ : Odrv4
    port map (
            O => \N__47337\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11\
        );

    \I__10509\ : InMux
    port map (
            O => \N__47334\,
            I => \N__47330\
        );

    \I__10508\ : InMux
    port map (
            O => \N__47333\,
            I => \N__47327\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__47330\,
            I => \N__47322\
        );

    \I__10506\ : LocalMux
    port map (
            O => \N__47327\,
            I => \N__47322\
        );

    \I__10505\ : Span4Mux_h
    port map (
            O => \N__47322\,
            I => \N__47319\
        );

    \I__10504\ : Odrv4
    port map (
            O => \N__47319\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49\
        );

    \I__10503\ : InMux
    port map (
            O => \N__47316\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10\
        );

    \I__10502\ : InMux
    port map (
            O => \N__47313\,
            I => \N__47309\
        );

    \I__10501\ : InMux
    port map (
            O => \N__47312\,
            I => \N__47306\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__47309\,
            I => \N__47301\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__47306\,
            I => \N__47301\
        );

    \I__10498\ : Span4Mux_h
    port map (
            O => \N__47301\,
            I => \N__47298\
        );

    \I__10497\ : Odrv4
    port map (
            O => \N__47298\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59\
        );

    \I__10496\ : InMux
    port map (
            O => \N__47295\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11\
        );

    \I__10495\ : InMux
    port map (
            O => \N__47292\,
            I => \N__47288\
        );

    \I__10494\ : InMux
    port map (
            O => \N__47291\,
            I => \N__47285\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__47288\,
            I => \N__47282\
        );

    \I__10492\ : LocalMux
    port map (
            O => \N__47285\,
            I => \N__47279\
        );

    \I__10491\ : Span4Mux_v
    port map (
            O => \N__47282\,
            I => \N__47274\
        );

    \I__10490\ : Span4Mux_v
    port map (
            O => \N__47279\,
            I => \N__47274\
        );

    \I__10489\ : Odrv4
    port map (
            O => \N__47274\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69\
        );

    \I__10488\ : InMux
    port map (
            O => \N__47271\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12\
        );

    \I__10487\ : InMux
    port map (
            O => \N__47268\,
            I => \N__47265\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__47265\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14\
        );

    \I__10485\ : InMux
    port map (
            O => \N__47262\,
            I => \N__47258\
        );

    \I__10484\ : InMux
    port map (
            O => \N__47261\,
            I => \N__47255\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__47258\,
            I => \N__47250\
        );

    \I__10482\ : LocalMux
    port map (
            O => \N__47255\,
            I => \N__47250\
        );

    \I__10481\ : Span4Mux_h
    port map (
            O => \N__47250\,
            I => \N__47247\
        );

    \I__10480\ : Odrv4
    port map (
            O => \N__47247\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79\
        );

    \I__10479\ : InMux
    port map (
            O => \N__47244\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13\
        );

    \I__10478\ : InMux
    port map (
            O => \N__47241\,
            I => \N__47238\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__47238\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15\
        );

    \I__10476\ : InMux
    port map (
            O => \N__47235\,
            I => \N__47231\
        );

    \I__10475\ : InMux
    port map (
            O => \N__47234\,
            I => \N__47228\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__47231\,
            I => \N__47223\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__47228\,
            I => \N__47223\
        );

    \I__10472\ : Odrv12
    port map (
            O => \N__47223\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099\
        );

    \I__10471\ : InMux
    port map (
            O => \N__47220\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14\
        );

    \I__10470\ : InMux
    port map (
            O => \N__47217\,
            I => \N__47214\
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__47214\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16\
        );

    \I__10468\ : InMux
    port map (
            O => \N__47211\,
            I => \N__47207\
        );

    \I__10467\ : InMux
    port map (
            O => \N__47210\,
            I => \N__47204\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__47207\,
            I => \N__47199\
        );

    \I__10465\ : LocalMux
    port map (
            O => \N__47204\,
            I => \N__47199\
        );

    \I__10464\ : Span4Mux_h
    port map (
            O => \N__47199\,
            I => \N__47196\
        );

    \I__10463\ : Span4Mux_v
    port map (
            O => \N__47196\,
            I => \N__47193\
        );

    \I__10462\ : Odrv4
    port map (
            O => \N__47193\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9\
        );

    \I__10461\ : InMux
    port map (
            O => \N__47190\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15\
        );

    \I__10460\ : InMux
    port map (
            O => \N__47187\,
            I => \N__47184\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__47184\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17\
        );

    \I__10458\ : InMux
    port map (
            O => \N__47181\,
            I => \N__47177\
        );

    \I__10457\ : InMux
    port map (
            O => \N__47180\,
            I => \N__47174\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__47177\,
            I => \N__47169\
        );

    \I__10455\ : LocalMux
    port map (
            O => \N__47174\,
            I => \N__47169\
        );

    \I__10454\ : Odrv12
    port map (
            O => \N__47169\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9\
        );

    \I__10453\ : InMux
    port map (
            O => \N__47166\,
            I => \bfn_17_14_0_\
        );

    \I__10452\ : InMux
    port map (
            O => \N__47163\,
            I => \N__47160\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__47160\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3\
        );

    \I__10450\ : InMux
    port map (
            O => \N__47157\,
            I => \N__47154\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__47154\,
            I => \N__47150\
        );

    \I__10448\ : CascadeMux
    port map (
            O => \N__47153\,
            I => \N__47146\
        );

    \I__10447\ : Span4Mux_v
    port map (
            O => \N__47150\,
            I => \N__47143\
        );

    \I__10446\ : InMux
    port map (
            O => \N__47149\,
            I => \N__47140\
        );

    \I__10445\ : InMux
    port map (
            O => \N__47146\,
            I => \N__47137\
        );

    \I__10444\ : Span4Mux_h
    port map (
            O => \N__47143\,
            I => \N__47134\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__47140\,
            I => \N__47131\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__47137\,
            I => \N__47128\
        );

    \I__10441\ : Span4Mux_h
    port map (
            O => \N__47134\,
            I => \N__47125\
        );

    \I__10440\ : Span4Mux_h
    port map (
            O => \N__47131\,
            I => \N__47120\
        );

    \I__10439\ : Span4Mux_h
    port map (
            O => \N__47128\,
            I => \N__47120\
        );

    \I__10438\ : Odrv4
    port map (
            O => \N__47125\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\
        );

    \I__10437\ : Odrv4
    port map (
            O => \N__47120\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\
        );

    \I__10436\ : InMux
    port map (
            O => \N__47115\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2\
        );

    \I__10435\ : InMux
    port map (
            O => \N__47112\,
            I => \N__47109\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__47109\,
            I => \N__47106\
        );

    \I__10433\ : Odrv4
    port map (
            O => \N__47106\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4\
        );

    \I__10432\ : InMux
    port map (
            O => \N__47103\,
            I => \N__47099\
        );

    \I__10431\ : InMux
    port map (
            O => \N__47102\,
            I => \N__47096\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__47099\,
            I => \N__47091\
        );

    \I__10429\ : LocalMux
    port map (
            O => \N__47096\,
            I => \N__47091\
        );

    \I__10428\ : Span4Mux_v
    port map (
            O => \N__47091\,
            I => \N__47088\
        );

    \I__10427\ : Odrv4
    port map (
            O => \N__47088\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0\
        );

    \I__10426\ : InMux
    port map (
            O => \N__47085\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3\
        );

    \I__10425\ : InMux
    port map (
            O => \N__47082\,
            I => \N__47078\
        );

    \I__10424\ : InMux
    port map (
            O => \N__47081\,
            I => \N__47075\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__47078\,
            I => \N__47070\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__47075\,
            I => \N__47070\
        );

    \I__10421\ : Odrv12
    port map (
            O => \N__47070\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0\
        );

    \I__10420\ : InMux
    port map (
            O => \N__47067\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4\
        );

    \I__10419\ : InMux
    port map (
            O => \N__47064\,
            I => \N__47061\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__47061\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6\
        );

    \I__10417\ : InMux
    port map (
            O => \N__47058\,
            I => \N__47054\
        );

    \I__10416\ : InMux
    port map (
            O => \N__47057\,
            I => \N__47051\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__47054\,
            I => \N__47046\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__47051\,
            I => \N__47046\
        );

    \I__10413\ : Odrv12
    port map (
            O => \N__47046\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0\
        );

    \I__10412\ : InMux
    port map (
            O => \N__47043\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5\
        );

    \I__10411\ : InMux
    port map (
            O => \N__47040\,
            I => \N__47037\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__47037\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7\
        );

    \I__10409\ : InMux
    port map (
            O => \N__47034\,
            I => \N__47030\
        );

    \I__10408\ : InMux
    port map (
            O => \N__47033\,
            I => \N__47027\
        );

    \I__10407\ : LocalMux
    port map (
            O => \N__47030\,
            I => \N__47022\
        );

    \I__10406\ : LocalMux
    port map (
            O => \N__47027\,
            I => \N__47022\
        );

    \I__10405\ : Span4Mux_v
    port map (
            O => \N__47022\,
            I => \N__47019\
        );

    \I__10404\ : Odrv4
    port map (
            O => \N__47019\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26\
        );

    \I__10403\ : InMux
    port map (
            O => \N__47016\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6\
        );

    \I__10402\ : InMux
    port map (
            O => \N__47013\,
            I => \N__47010\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__47010\,
            I => \N__47007\
        );

    \I__10400\ : Span4Mux_h
    port map (
            O => \N__47007\,
            I => \N__47004\
        );

    \I__10399\ : Odrv4
    port map (
            O => \N__47004\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8\
        );

    \I__10398\ : InMux
    port map (
            O => \N__47001\,
            I => \N__46997\
        );

    \I__10397\ : InMux
    port map (
            O => \N__47000\,
            I => \N__46994\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__46997\,
            I => \N__46989\
        );

    \I__10395\ : LocalMux
    port map (
            O => \N__46994\,
            I => \N__46989\
        );

    \I__10394\ : Span4Mux_v
    port map (
            O => \N__46989\,
            I => \N__46986\
        );

    \I__10393\ : Odrv4
    port map (
            O => \N__46986\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381\
        );

    \I__10392\ : InMux
    port map (
            O => \N__46983\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7\
        );

    \I__10391\ : InMux
    port map (
            O => \N__46980\,
            I => \N__46977\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__46977\,
            I => \N__46974\
        );

    \I__10389\ : Span4Mux_v
    port map (
            O => \N__46974\,
            I => \N__46971\
        );

    \I__10388\ : Odrv4
    port map (
            O => \N__46971\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9\
        );

    \I__10387\ : InMux
    port map (
            O => \N__46968\,
            I => \N__46964\
        );

    \I__10386\ : InMux
    port map (
            O => \N__46967\,
            I => \N__46961\
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__46964\,
            I => \N__46956\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__46961\,
            I => \N__46956\
        );

    \I__10383\ : Odrv12
    port map (
            O => \N__46956\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2\
        );

    \I__10382\ : InMux
    port map (
            O => \N__46953\,
            I => \bfn_17_13_0_\
        );

    \I__10381\ : InMux
    port map (
            O => \N__46950\,
            I => \N__46947\
        );

    \I__10380\ : LocalMux
    port map (
            O => \N__46947\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10\
        );

    \I__10379\ : InMux
    port map (
            O => \N__46944\,
            I => \N__46941\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__46941\,
            I => \N__46937\
        );

    \I__10377\ : InMux
    port map (
            O => \N__46940\,
            I => \N__46934\
        );

    \I__10376\ : Span4Mux_v
    port map (
            O => \N__46937\,
            I => \N__46929\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__46934\,
            I => \N__46929\
        );

    \I__10374\ : Odrv4
    port map (
            O => \N__46929\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_22
        );

    \I__10373\ : InMux
    port map (
            O => \N__46926\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21\
        );

    \I__10372\ : InMux
    port map (
            O => \N__46923\,
            I => \N__46919\
        );

    \I__10371\ : InMux
    port map (
            O => \N__46922\,
            I => \N__46916\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__46919\,
            I => \N__46913\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__46916\,
            I => \N__46910\
        );

    \I__10368\ : Span4Mux_h
    port map (
            O => \N__46913\,
            I => \N__46907\
        );

    \I__10367\ : Span4Mux_h
    port map (
            O => \N__46910\,
            I => \N__46904\
        );

    \I__10366\ : Odrv4
    port map (
            O => \N__46907\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_23
        );

    \I__10365\ : Odrv4
    port map (
            O => \N__46904\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_23
        );

    \I__10364\ : InMux
    port map (
            O => \N__46899\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22\
        );

    \I__10363\ : InMux
    port map (
            O => \N__46896\,
            I => \bfn_17_11_0_\
        );

    \I__10362\ : InMux
    port map (
            O => \N__46893\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24\
        );

    \I__10361\ : InMux
    port map (
            O => \N__46890\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25\
        );

    \I__10360\ : CascadeMux
    port map (
            O => \N__46887\,
            I => \N__46869\
        );

    \I__10359\ : CascadeMux
    port map (
            O => \N__46886\,
            I => \N__46866\
        );

    \I__10358\ : CascadeMux
    port map (
            O => \N__46885\,
            I => \N__46863\
        );

    \I__10357\ : CascadeMux
    port map (
            O => \N__46884\,
            I => \N__46860\
        );

    \I__10356\ : CascadeMux
    port map (
            O => \N__46883\,
            I => \N__46857\
        );

    \I__10355\ : CascadeMux
    port map (
            O => \N__46882\,
            I => \N__46854\
        );

    \I__10354\ : CascadeMux
    port map (
            O => \N__46881\,
            I => \N__46833\
        );

    \I__10353\ : CascadeMux
    port map (
            O => \N__46880\,
            I => \N__46830\
        );

    \I__10352\ : CascadeMux
    port map (
            O => \N__46879\,
            I => \N__46825\
        );

    \I__10351\ : CascadeMux
    port map (
            O => \N__46878\,
            I => \N__46822\
        );

    \I__10350\ : CascadeMux
    port map (
            O => \N__46877\,
            I => \N__46819\
        );

    \I__10349\ : CascadeMux
    port map (
            O => \N__46876\,
            I => \N__46816\
        );

    \I__10348\ : CascadeMux
    port map (
            O => \N__46875\,
            I => \N__46813\
        );

    \I__10347\ : CascadeMux
    port map (
            O => \N__46874\,
            I => \N__46810\
        );

    \I__10346\ : CascadeMux
    port map (
            O => \N__46873\,
            I => \N__46807\
        );

    \I__10345\ : CascadeMux
    port map (
            O => \N__46872\,
            I => \N__46804\
        );

    \I__10344\ : InMux
    port map (
            O => \N__46869\,
            I => \N__46799\
        );

    \I__10343\ : InMux
    port map (
            O => \N__46866\,
            I => \N__46799\
        );

    \I__10342\ : InMux
    port map (
            O => \N__46863\,
            I => \N__46790\
        );

    \I__10341\ : InMux
    port map (
            O => \N__46860\,
            I => \N__46790\
        );

    \I__10340\ : InMux
    port map (
            O => \N__46857\,
            I => \N__46790\
        );

    \I__10339\ : InMux
    port map (
            O => \N__46854\,
            I => \N__46790\
        );

    \I__10338\ : CascadeMux
    port map (
            O => \N__46853\,
            I => \N__46787\
        );

    \I__10337\ : CascadeMux
    port map (
            O => \N__46852\,
            I => \N__46784\
        );

    \I__10336\ : CascadeMux
    port map (
            O => \N__46851\,
            I => \N__46781\
        );

    \I__10335\ : CascadeMux
    port map (
            O => \N__46850\,
            I => \N__46778\
        );

    \I__10334\ : CascadeMux
    port map (
            O => \N__46849\,
            I => \N__46775\
        );

    \I__10333\ : CascadeMux
    port map (
            O => \N__46848\,
            I => \N__46772\
        );

    \I__10332\ : CascadeMux
    port map (
            O => \N__46847\,
            I => \N__46754\
        );

    \I__10331\ : CascadeMux
    port map (
            O => \N__46846\,
            I => \N__46751\
        );

    \I__10330\ : CascadeMux
    port map (
            O => \N__46845\,
            I => \N__46748\
        );

    \I__10329\ : CascadeMux
    port map (
            O => \N__46844\,
            I => \N__46745\
        );

    \I__10328\ : CascadeMux
    port map (
            O => \N__46843\,
            I => \N__46742\
        );

    \I__10327\ : CascadeMux
    port map (
            O => \N__46842\,
            I => \N__46739\
        );

    \I__10326\ : CascadeMux
    port map (
            O => \N__46841\,
            I => \N__46736\
        );

    \I__10325\ : CascadeMux
    port map (
            O => \N__46840\,
            I => \N__46733\
        );

    \I__10324\ : CascadeMux
    port map (
            O => \N__46839\,
            I => \N__46730\
        );

    \I__10323\ : CascadeMux
    port map (
            O => \N__46838\,
            I => \N__46727\
        );

    \I__10322\ : CascadeMux
    port map (
            O => \N__46837\,
            I => \N__46724\
        );

    \I__10321\ : CascadeMux
    port map (
            O => \N__46836\,
            I => \N__46721\
        );

    \I__10320\ : InMux
    port map (
            O => \N__46833\,
            I => \N__46718\
        );

    \I__10319\ : InMux
    port map (
            O => \N__46830\,
            I => \N__46713\
        );

    \I__10318\ : InMux
    port map (
            O => \N__46829\,
            I => \N__46713\
        );

    \I__10317\ : InMux
    port map (
            O => \N__46828\,
            I => \N__46710\
        );

    \I__10316\ : InMux
    port map (
            O => \N__46825\,
            I => \N__46705\
        );

    \I__10315\ : InMux
    port map (
            O => \N__46822\,
            I => \N__46705\
        );

    \I__10314\ : InMux
    port map (
            O => \N__46819\,
            I => \N__46700\
        );

    \I__10313\ : InMux
    port map (
            O => \N__46816\,
            I => \N__46700\
        );

    \I__10312\ : InMux
    port map (
            O => \N__46813\,
            I => \N__46691\
        );

    \I__10311\ : InMux
    port map (
            O => \N__46810\,
            I => \N__46691\
        );

    \I__10310\ : InMux
    port map (
            O => \N__46807\,
            I => \N__46691\
        );

    \I__10309\ : InMux
    port map (
            O => \N__46804\,
            I => \N__46691\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__46799\,
            I => \N__46681\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__46790\,
            I => \N__46678\
        );

    \I__10306\ : InMux
    port map (
            O => \N__46787\,
            I => \N__46669\
        );

    \I__10305\ : InMux
    port map (
            O => \N__46784\,
            I => \N__46669\
        );

    \I__10304\ : InMux
    port map (
            O => \N__46781\,
            I => \N__46669\
        );

    \I__10303\ : InMux
    port map (
            O => \N__46778\,
            I => \N__46669\
        );

    \I__10302\ : InMux
    port map (
            O => \N__46775\,
            I => \N__46664\
        );

    \I__10301\ : InMux
    port map (
            O => \N__46772\,
            I => \N__46664\
        );

    \I__10300\ : CascadeMux
    port map (
            O => \N__46771\,
            I => \N__46661\
        );

    \I__10299\ : CascadeMux
    port map (
            O => \N__46770\,
            I => \N__46658\
        );

    \I__10298\ : CascadeMux
    port map (
            O => \N__46769\,
            I => \N__46655\
        );

    \I__10297\ : CascadeMux
    port map (
            O => \N__46768\,
            I => \N__46652\
        );

    \I__10296\ : CascadeMux
    port map (
            O => \N__46767\,
            I => \N__46649\
        );

    \I__10295\ : CascadeMux
    port map (
            O => \N__46766\,
            I => \N__46646\
        );

    \I__10294\ : CascadeMux
    port map (
            O => \N__46765\,
            I => \N__46643\
        );

    \I__10293\ : CascadeMux
    port map (
            O => \N__46764\,
            I => \N__46640\
        );

    \I__10292\ : CascadeMux
    port map (
            O => \N__46763\,
            I => \N__46637\
        );

    \I__10291\ : CascadeMux
    port map (
            O => \N__46762\,
            I => \N__46634\
        );

    \I__10290\ : CascadeMux
    port map (
            O => \N__46761\,
            I => \N__46631\
        );

    \I__10289\ : CascadeMux
    port map (
            O => \N__46760\,
            I => \N__46628\
        );

    \I__10288\ : CascadeMux
    port map (
            O => \N__46759\,
            I => \N__46625\
        );

    \I__10287\ : CascadeMux
    port map (
            O => \N__46758\,
            I => \N__46622\
        );

    \I__10286\ : CascadeMux
    port map (
            O => \N__46757\,
            I => \N__46619\
        );

    \I__10285\ : InMux
    port map (
            O => \N__46754\,
            I => \N__46610\
        );

    \I__10284\ : InMux
    port map (
            O => \N__46751\,
            I => \N__46610\
        );

    \I__10283\ : InMux
    port map (
            O => \N__46748\,
            I => \N__46610\
        );

    \I__10282\ : InMux
    port map (
            O => \N__46745\,
            I => \N__46610\
        );

    \I__10281\ : InMux
    port map (
            O => \N__46742\,
            I => \N__46601\
        );

    \I__10280\ : InMux
    port map (
            O => \N__46739\,
            I => \N__46601\
        );

    \I__10279\ : InMux
    port map (
            O => \N__46736\,
            I => \N__46601\
        );

    \I__10278\ : InMux
    port map (
            O => \N__46733\,
            I => \N__46601\
        );

    \I__10277\ : InMux
    port map (
            O => \N__46730\,
            I => \N__46592\
        );

    \I__10276\ : InMux
    port map (
            O => \N__46727\,
            I => \N__46592\
        );

    \I__10275\ : InMux
    port map (
            O => \N__46724\,
            I => \N__46592\
        );

    \I__10274\ : InMux
    port map (
            O => \N__46721\,
            I => \N__46592\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__46718\,
            I => \N__46587\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__46713\,
            I => \N__46587\
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__46710\,
            I => \N__46573\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__46705\,
            I => \N__46566\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__46700\,
            I => \N__46566\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__46691\,
            I => \N__46566\
        );

    \I__10267\ : CascadeMux
    port map (
            O => \N__46690\,
            I => \N__46563\
        );

    \I__10266\ : CascadeMux
    port map (
            O => \N__46689\,
            I => \N__46560\
        );

    \I__10265\ : CascadeMux
    port map (
            O => \N__46688\,
            I => \N__46557\
        );

    \I__10264\ : CascadeMux
    port map (
            O => \N__46687\,
            I => \N__46554\
        );

    \I__10263\ : CascadeMux
    port map (
            O => \N__46686\,
            I => \N__46551\
        );

    \I__10262\ : CascadeMux
    port map (
            O => \N__46685\,
            I => \N__46548\
        );

    \I__10261\ : CascadeMux
    port map (
            O => \N__46684\,
            I => \N__46545\
        );

    \I__10260\ : Span4Mux_v
    port map (
            O => \N__46681\,
            I => \N__46538\
        );

    \I__10259\ : Span4Mux_h
    port map (
            O => \N__46678\,
            I => \N__46538\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__46669\,
            I => \N__46538\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__46664\,
            I => \N__46535\
        );

    \I__10256\ : InMux
    port map (
            O => \N__46661\,
            I => \N__46526\
        );

    \I__10255\ : InMux
    port map (
            O => \N__46658\,
            I => \N__46526\
        );

    \I__10254\ : InMux
    port map (
            O => \N__46655\,
            I => \N__46526\
        );

    \I__10253\ : InMux
    port map (
            O => \N__46652\,
            I => \N__46526\
        );

    \I__10252\ : InMux
    port map (
            O => \N__46649\,
            I => \N__46517\
        );

    \I__10251\ : InMux
    port map (
            O => \N__46646\,
            I => \N__46517\
        );

    \I__10250\ : InMux
    port map (
            O => \N__46643\,
            I => \N__46517\
        );

    \I__10249\ : InMux
    port map (
            O => \N__46640\,
            I => \N__46517\
        );

    \I__10248\ : InMux
    port map (
            O => \N__46637\,
            I => \N__46510\
        );

    \I__10247\ : InMux
    port map (
            O => \N__46634\,
            I => \N__46510\
        );

    \I__10246\ : InMux
    port map (
            O => \N__46631\,
            I => \N__46510\
        );

    \I__10245\ : InMux
    port map (
            O => \N__46628\,
            I => \N__46501\
        );

    \I__10244\ : InMux
    port map (
            O => \N__46625\,
            I => \N__46501\
        );

    \I__10243\ : InMux
    port map (
            O => \N__46622\,
            I => \N__46501\
        );

    \I__10242\ : InMux
    port map (
            O => \N__46619\,
            I => \N__46501\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__46610\,
            I => \N__46494\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__46601\,
            I => \N__46494\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__46592\,
            I => \N__46494\
        );

    \I__10238\ : Span4Mux_v
    port map (
            O => \N__46587\,
            I => \N__46491\
        );

    \I__10237\ : InMux
    port map (
            O => \N__46586\,
            I => \N__46475\
        );

    \I__10236\ : InMux
    port map (
            O => \N__46585\,
            I => \N__46468\
        );

    \I__10235\ : InMux
    port map (
            O => \N__46584\,
            I => \N__46468\
        );

    \I__10234\ : InMux
    port map (
            O => \N__46583\,
            I => \N__46468\
        );

    \I__10233\ : InMux
    port map (
            O => \N__46582\,
            I => \N__46459\
        );

    \I__10232\ : InMux
    port map (
            O => \N__46581\,
            I => \N__46459\
        );

    \I__10231\ : InMux
    port map (
            O => \N__46580\,
            I => \N__46459\
        );

    \I__10230\ : InMux
    port map (
            O => \N__46579\,
            I => \N__46459\
        );

    \I__10229\ : InMux
    port map (
            O => \N__46578\,
            I => \N__46456\
        );

    \I__10228\ : InMux
    port map (
            O => \N__46577\,
            I => \N__46453\
        );

    \I__10227\ : InMux
    port map (
            O => \N__46576\,
            I => \N__46450\
        );

    \I__10226\ : Span12Mux_s11_v
    port map (
            O => \N__46573\,
            I => \N__46439\
        );

    \I__10225\ : Span4Mux_v
    port map (
            O => \N__46566\,
            I => \N__46436\
        );

    \I__10224\ : InMux
    port map (
            O => \N__46563\,
            I => \N__46429\
        );

    \I__10223\ : InMux
    port map (
            O => \N__46560\,
            I => \N__46429\
        );

    \I__10222\ : InMux
    port map (
            O => \N__46557\,
            I => \N__46429\
        );

    \I__10221\ : InMux
    port map (
            O => \N__46554\,
            I => \N__46420\
        );

    \I__10220\ : InMux
    port map (
            O => \N__46551\,
            I => \N__46420\
        );

    \I__10219\ : InMux
    port map (
            O => \N__46548\,
            I => \N__46420\
        );

    \I__10218\ : InMux
    port map (
            O => \N__46545\,
            I => \N__46420\
        );

    \I__10217\ : Span4Mux_v
    port map (
            O => \N__46538\,
            I => \N__46417\
        );

    \I__10216\ : Span4Mux_v
    port map (
            O => \N__46535\,
            I => \N__46412\
        );

    \I__10215\ : LocalMux
    port map (
            O => \N__46526\,
            I => \N__46412\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__46517\,
            I => \N__46405\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__46510\,
            I => \N__46405\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__46501\,
            I => \N__46405\
        );

    \I__10211\ : Span4Mux_v
    port map (
            O => \N__46494\,
            I => \N__46402\
        );

    \I__10210\ : Sp12to4
    port map (
            O => \N__46491\,
            I => \N__46399\
        );

    \I__10209\ : InMux
    port map (
            O => \N__46490\,
            I => \N__46394\
        );

    \I__10208\ : InMux
    port map (
            O => \N__46489\,
            I => \N__46394\
        );

    \I__10207\ : CascadeMux
    port map (
            O => \N__46488\,
            I => \N__46390\
        );

    \I__10206\ : CascadeMux
    port map (
            O => \N__46487\,
            I => \N__46386\
        );

    \I__10205\ : CascadeMux
    port map (
            O => \N__46486\,
            I => \N__46382\
        );

    \I__10204\ : CascadeMux
    port map (
            O => \N__46485\,
            I => \N__46377\
        );

    \I__10203\ : CascadeMux
    port map (
            O => \N__46484\,
            I => \N__46373\
        );

    \I__10202\ : CascadeMux
    port map (
            O => \N__46483\,
            I => \N__46369\
        );

    \I__10201\ : CascadeMux
    port map (
            O => \N__46482\,
            I => \N__46365\
        );

    \I__10200\ : CascadeMux
    port map (
            O => \N__46481\,
            I => \N__46362\
        );

    \I__10199\ : CascadeMux
    port map (
            O => \N__46480\,
            I => \N__46358\
        );

    \I__10198\ : CascadeMux
    port map (
            O => \N__46479\,
            I => \N__46354\
        );

    \I__10197\ : CascadeMux
    port map (
            O => \N__46478\,
            I => \N__46350\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__46475\,
            I => \N__46335\
        );

    \I__10195\ : LocalMux
    port map (
            O => \N__46468\,
            I => \N__46335\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__46459\,
            I => \N__46335\
        );

    \I__10193\ : LocalMux
    port map (
            O => \N__46456\,
            I => \N__46330\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__46453\,
            I => \N__46330\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__46450\,
            I => \N__46327\
        );

    \I__10190\ : InMux
    port map (
            O => \N__46449\,
            I => \N__46324\
        );

    \I__10189\ : InMux
    port map (
            O => \N__46448\,
            I => \N__46317\
        );

    \I__10188\ : InMux
    port map (
            O => \N__46447\,
            I => \N__46317\
        );

    \I__10187\ : InMux
    port map (
            O => \N__46446\,
            I => \N__46317\
        );

    \I__10186\ : InMux
    port map (
            O => \N__46445\,
            I => \N__46308\
        );

    \I__10185\ : InMux
    port map (
            O => \N__46444\,
            I => \N__46308\
        );

    \I__10184\ : InMux
    port map (
            O => \N__46443\,
            I => \N__46308\
        );

    \I__10183\ : InMux
    port map (
            O => \N__46442\,
            I => \N__46308\
        );

    \I__10182\ : Span12Mux_v
    port map (
            O => \N__46439\,
            I => \N__46301\
        );

    \I__10181\ : Sp12to4
    port map (
            O => \N__46436\,
            I => \N__46294\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__46429\,
            I => \N__46294\
        );

    \I__10179\ : LocalMux
    port map (
            O => \N__46420\,
            I => \N__46294\
        );

    \I__10178\ : Span4Mux_h
    port map (
            O => \N__46417\,
            I => \N__46289\
        );

    \I__10177\ : Span4Mux_v
    port map (
            O => \N__46412\,
            I => \N__46289\
        );

    \I__10176\ : Span4Mux_v
    port map (
            O => \N__46405\,
            I => \N__46286\
        );

    \I__10175\ : Sp12to4
    port map (
            O => \N__46402\,
            I => \N__46283\
        );

    \I__10174\ : Span12Mux_h
    port map (
            O => \N__46399\,
            I => \N__46278\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__46394\,
            I => \N__46278\
        );

    \I__10172\ : InMux
    port map (
            O => \N__46393\,
            I => \N__46263\
        );

    \I__10171\ : InMux
    port map (
            O => \N__46390\,
            I => \N__46263\
        );

    \I__10170\ : InMux
    port map (
            O => \N__46389\,
            I => \N__46263\
        );

    \I__10169\ : InMux
    port map (
            O => \N__46386\,
            I => \N__46263\
        );

    \I__10168\ : InMux
    port map (
            O => \N__46385\,
            I => \N__46263\
        );

    \I__10167\ : InMux
    port map (
            O => \N__46382\,
            I => \N__46263\
        );

    \I__10166\ : InMux
    port map (
            O => \N__46381\,
            I => \N__46263\
        );

    \I__10165\ : InMux
    port map (
            O => \N__46380\,
            I => \N__46246\
        );

    \I__10164\ : InMux
    port map (
            O => \N__46377\,
            I => \N__46246\
        );

    \I__10163\ : InMux
    port map (
            O => \N__46376\,
            I => \N__46246\
        );

    \I__10162\ : InMux
    port map (
            O => \N__46373\,
            I => \N__46246\
        );

    \I__10161\ : InMux
    port map (
            O => \N__46372\,
            I => \N__46246\
        );

    \I__10160\ : InMux
    port map (
            O => \N__46369\,
            I => \N__46246\
        );

    \I__10159\ : InMux
    port map (
            O => \N__46368\,
            I => \N__46246\
        );

    \I__10158\ : InMux
    port map (
            O => \N__46365\,
            I => \N__46246\
        );

    \I__10157\ : InMux
    port map (
            O => \N__46362\,
            I => \N__46229\
        );

    \I__10156\ : InMux
    port map (
            O => \N__46361\,
            I => \N__46229\
        );

    \I__10155\ : InMux
    port map (
            O => \N__46358\,
            I => \N__46229\
        );

    \I__10154\ : InMux
    port map (
            O => \N__46357\,
            I => \N__46229\
        );

    \I__10153\ : InMux
    port map (
            O => \N__46354\,
            I => \N__46229\
        );

    \I__10152\ : InMux
    port map (
            O => \N__46353\,
            I => \N__46229\
        );

    \I__10151\ : InMux
    port map (
            O => \N__46350\,
            I => \N__46229\
        );

    \I__10150\ : InMux
    port map (
            O => \N__46349\,
            I => \N__46229\
        );

    \I__10149\ : InMux
    port map (
            O => \N__46348\,
            I => \N__46222\
        );

    \I__10148\ : InMux
    port map (
            O => \N__46347\,
            I => \N__46222\
        );

    \I__10147\ : InMux
    port map (
            O => \N__46346\,
            I => \N__46222\
        );

    \I__10146\ : InMux
    port map (
            O => \N__46345\,
            I => \N__46213\
        );

    \I__10145\ : InMux
    port map (
            O => \N__46344\,
            I => \N__46213\
        );

    \I__10144\ : InMux
    port map (
            O => \N__46343\,
            I => \N__46213\
        );

    \I__10143\ : InMux
    port map (
            O => \N__46342\,
            I => \N__46213\
        );

    \I__10142\ : Span12Mux_v
    port map (
            O => \N__46335\,
            I => \N__46210\
        );

    \I__10141\ : Span4Mux_v
    port map (
            O => \N__46330\,
            I => \N__46201\
        );

    \I__10140\ : Span4Mux_v
    port map (
            O => \N__46327\,
            I => \N__46201\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__46324\,
            I => \N__46201\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__46317\,
            I => \N__46201\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__46308\,
            I => \N__46198\
        );

    \I__10136\ : InMux
    port map (
            O => \N__46307\,
            I => \N__46193\
        );

    \I__10135\ : InMux
    port map (
            O => \N__46306\,
            I => \N__46193\
        );

    \I__10134\ : InMux
    port map (
            O => \N__46305\,
            I => \N__46190\
        );

    \I__10133\ : InMux
    port map (
            O => \N__46304\,
            I => \N__46187\
        );

    \I__10132\ : Span12Mux_h
    port map (
            O => \N__46301\,
            I => \N__46182\
        );

    \I__10131\ : Span12Mux_v
    port map (
            O => \N__46294\,
            I => \N__46182\
        );

    \I__10130\ : Sp12to4
    port map (
            O => \N__46289\,
            I => \N__46177\
        );

    \I__10129\ : Sp12to4
    port map (
            O => \N__46286\,
            I => \N__46177\
        );

    \I__10128\ : Span12Mux_h
    port map (
            O => \N__46283\,
            I => \N__46162\
        );

    \I__10127\ : Span12Mux_v
    port map (
            O => \N__46278\,
            I => \N__46162\
        );

    \I__10126\ : LocalMux
    port map (
            O => \N__46263\,
            I => \N__46162\
        );

    \I__10125\ : LocalMux
    port map (
            O => \N__46246\,
            I => \N__46162\
        );

    \I__10124\ : LocalMux
    port map (
            O => \N__46229\,
            I => \N__46162\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__46222\,
            I => \N__46162\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__46213\,
            I => \N__46162\
        );

    \I__10121\ : Span12Mux_h
    port map (
            O => \N__46210\,
            I => \N__46159\
        );

    \I__10120\ : Sp12to4
    port map (
            O => \N__46201\,
            I => \N__46154\
        );

    \I__10119\ : Sp12to4
    port map (
            O => \N__46198\,
            I => \N__46154\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__46193\,
            I => \N__46151\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__46190\,
            I => \N__46146\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__46187\,
            I => \N__46146\
        );

    \I__10115\ : Span12Mux_h
    port map (
            O => \N__46182\,
            I => \N__46139\
        );

    \I__10114\ : Span12Mux_h
    port map (
            O => \N__46177\,
            I => \N__46134\
        );

    \I__10113\ : Span12Mux_v
    port map (
            O => \N__46162\,
            I => \N__46134\
        );

    \I__10112\ : Span12Mux_h
    port map (
            O => \N__46159\,
            I => \N__46125\
        );

    \I__10111\ : Span12Mux_v
    port map (
            O => \N__46154\,
            I => \N__46125\
        );

    \I__10110\ : Sp12to4
    port map (
            O => \N__46151\,
            I => \N__46125\
        );

    \I__10109\ : Sp12to4
    port map (
            O => \N__46146\,
            I => \N__46125\
        );

    \I__10108\ : InMux
    port map (
            O => \N__46145\,
            I => \N__46122\
        );

    \I__10107\ : InMux
    port map (
            O => \N__46144\,
            I => \N__46117\
        );

    \I__10106\ : InMux
    port map (
            O => \N__46143\,
            I => \N__46117\
        );

    \I__10105\ : InMux
    port map (
            O => \N__46142\,
            I => \N__46114\
        );

    \I__10104\ : Odrv12
    port map (
            O => \N__46139\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10103\ : Odrv12
    port map (
            O => \N__46134\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10102\ : Odrv12
    port map (
            O => \N__46125\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__46122\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__46117\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__46114\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10098\ : InMux
    port map (
            O => \N__46101\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26\
        );

    \I__10097\ : InMux
    port map (
            O => \N__46098\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27\
        );

    \I__10096\ : InMux
    port map (
            O => \N__46095\,
            I => \N__46091\
        );

    \I__10095\ : InMux
    port map (
            O => \N__46094\,
            I => \N__46088\
        );

    \I__10094\ : LocalMux
    port map (
            O => \N__46091\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__46088\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10092\ : CascadeMux
    port map (
            O => \N__46083\,
            I => \N__46080\
        );

    \I__10091\ : InMux
    port map (
            O => \N__46080\,
            I => \N__46077\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__46077\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1\
        );

    \I__10089\ : InMux
    port map (
            O => \N__46074\,
            I => \N__46070\
        );

    \I__10088\ : InMux
    port map (
            O => \N__46073\,
            I => \N__46067\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__46070\,
            I => \N__46064\
        );

    \I__10086\ : LocalMux
    port map (
            O => \N__46067\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__10085\ : Odrv4
    port map (
            O => \N__46064\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__10084\ : InMux
    port map (
            O => \N__46059\,
            I => \N__46056\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__46056\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2\
        );

    \I__10082\ : InMux
    port map (
            O => \N__46053\,
            I => \N__46049\
        );

    \I__10081\ : InMux
    port map (
            O => \N__46052\,
            I => \N__46046\
        );

    \I__10080\ : LocalMux
    port map (
            O => \N__46049\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_13
        );

    \I__10079\ : LocalMux
    port map (
            O => \N__46046\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_13
        );

    \I__10078\ : InMux
    port map (
            O => \N__46041\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12\
        );

    \I__10077\ : InMux
    port map (
            O => \N__46038\,
            I => \N__46034\
        );

    \I__10076\ : InMux
    port map (
            O => \N__46037\,
            I => \N__46031\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__46034\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_14
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__46031\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_14
        );

    \I__10073\ : InMux
    port map (
            O => \N__46026\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13\
        );

    \I__10072\ : InMux
    port map (
            O => \N__46023\,
            I => \N__46019\
        );

    \I__10071\ : InMux
    port map (
            O => \N__46022\,
            I => \N__46016\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__46019\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_15
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__46016\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_15
        );

    \I__10068\ : InMux
    port map (
            O => \N__46011\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14\
        );

    \I__10067\ : InMux
    port map (
            O => \N__46008\,
            I => \bfn_17_10_0_\
        );

    \I__10066\ : InMux
    port map (
            O => \N__46005\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16\
        );

    \I__10065\ : InMux
    port map (
            O => \N__46002\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17\
        );

    \I__10064\ : InMux
    port map (
            O => \N__45999\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18\
        );

    \I__10063\ : InMux
    port map (
            O => \N__45996\,
            I => \N__45993\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__45993\,
            I => \N__45989\
        );

    \I__10061\ : InMux
    port map (
            O => \N__45992\,
            I => \N__45986\
        );

    \I__10060\ : Span4Mux_v
    port map (
            O => \N__45989\,
            I => \N__45981\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__45986\,
            I => \N__45981\
        );

    \I__10058\ : Odrv4
    port map (
            O => \N__45981\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_20
        );

    \I__10057\ : InMux
    port map (
            O => \N__45978\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19\
        );

    \I__10056\ : InMux
    port map (
            O => \N__45975\,
            I => \N__45971\
        );

    \I__10055\ : InMux
    port map (
            O => \N__45974\,
            I => \N__45968\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__45971\,
            I => \N__45965\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__45968\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_21
        );

    \I__10052\ : Odrv4
    port map (
            O => \N__45965\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_21
        );

    \I__10051\ : InMux
    port map (
            O => \N__45960\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20\
        );

    \I__10050\ : InMux
    port map (
            O => \N__45957\,
            I => \N__45954\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__45954\,
            I => \N__45950\
        );

    \I__10048\ : InMux
    port map (
            O => \N__45953\,
            I => \N__45947\
        );

    \I__10047\ : Odrv4
    port map (
            O => \N__45950\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_5
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__45947\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_5
        );

    \I__10045\ : InMux
    port map (
            O => \N__45942\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4\
        );

    \I__10044\ : InMux
    port map (
            O => \N__45939\,
            I => \N__45936\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__45936\,
            I => \N__45932\
        );

    \I__10042\ : InMux
    port map (
            O => \N__45935\,
            I => \N__45929\
        );

    \I__10041\ : Span4Mux_v
    port map (
            O => \N__45932\,
            I => \N__45924\
        );

    \I__10040\ : LocalMux
    port map (
            O => \N__45929\,
            I => \N__45924\
        );

    \I__10039\ : Odrv4
    port map (
            O => \N__45924\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_6
        );

    \I__10038\ : InMux
    port map (
            O => \N__45921\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5\
        );

    \I__10037\ : InMux
    port map (
            O => \N__45918\,
            I => \N__45915\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__45915\,
            I => \N__45911\
        );

    \I__10035\ : InMux
    port map (
            O => \N__45914\,
            I => \N__45908\
        );

    \I__10034\ : Odrv4
    port map (
            O => \N__45911\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_7
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__45908\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_7
        );

    \I__10032\ : InMux
    port map (
            O => \N__45903\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6\
        );

    \I__10031\ : InMux
    port map (
            O => \N__45900\,
            I => \N__45897\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__45897\,
            I => \N__45893\
        );

    \I__10029\ : InMux
    port map (
            O => \N__45896\,
            I => \N__45890\
        );

    \I__10028\ : Odrv4
    port map (
            O => \N__45893\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_8
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__45890\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_8
        );

    \I__10026\ : InMux
    port map (
            O => \N__45885\,
            I => \bfn_17_9_0_\
        );

    \I__10025\ : InMux
    port map (
            O => \N__45882\,
            I => \N__45878\
        );

    \I__10024\ : InMux
    port map (
            O => \N__45881\,
            I => \N__45875\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__45878\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_9
        );

    \I__10022\ : LocalMux
    port map (
            O => \N__45875\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_9
        );

    \I__10021\ : InMux
    port map (
            O => \N__45870\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8\
        );

    \I__10020\ : InMux
    port map (
            O => \N__45867\,
            I => \N__45863\
        );

    \I__10019\ : InMux
    port map (
            O => \N__45866\,
            I => \N__45860\
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__45863\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_10
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__45860\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_10
        );

    \I__10016\ : InMux
    port map (
            O => \N__45855\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9\
        );

    \I__10015\ : InMux
    port map (
            O => \N__45852\,
            I => \N__45848\
        );

    \I__10014\ : InMux
    port map (
            O => \N__45851\,
            I => \N__45845\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__45848\,
            I => \N__45842\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__45845\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_11
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__45842\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_11
        );

    \I__10010\ : InMux
    port map (
            O => \N__45837\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10\
        );

    \I__10009\ : InMux
    port map (
            O => \N__45834\,
            I => \N__45831\
        );

    \I__10008\ : LocalMux
    port map (
            O => \N__45831\,
            I => \N__45827\
        );

    \I__10007\ : InMux
    port map (
            O => \N__45830\,
            I => \N__45824\
        );

    \I__10006\ : Odrv4
    port map (
            O => \N__45827\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_12
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__45824\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_12
        );

    \I__10004\ : InMux
    port map (
            O => \N__45819\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11\
        );

    \I__10003\ : InMux
    port map (
            O => \N__45816\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14\
        );

    \I__10002\ : InMux
    port map (
            O => \N__45813\,
            I => \N__45810\
        );

    \I__10001\ : LocalMux
    port map (
            O => \N__45810\,
            I => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\
        );

    \I__10000\ : InMux
    port map (
            O => \N__45807\,
            I => \N__45804\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__45804\,
            I => \N__45801\
        );

    \I__9998\ : Odrv12
    port map (
            O => \N__45801\,
            I => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\
        );

    \I__9997\ : InMux
    port map (
            O => \N__45798\,
            I => \bfn_16_30_0_\
        );

    \I__9996\ : IoInMux
    port map (
            O => \N__45795\,
            I => \N__45792\
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__45792\,
            I => \GB_BUFFER_red_c_g_THRU_CO\
        );

    \I__9994\ : InMux
    port map (
            O => \N__45789\,
            I => \N__45783\
        );

    \I__9993\ : InMux
    port map (
            O => \N__45788\,
            I => \N__45783\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__45783\,
            I => \N__45780\
        );

    \I__9991\ : Span4Mux_h
    port map (
            O => \N__45780\,
            I => \N__45777\
        );

    \I__9990\ : Odrv4
    port map (
            O => \N__45777\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_23\
        );

    \I__9989\ : InMux
    port map (
            O => \N__45774\,
            I => \N__45771\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__45771\,
            I => \phase_controller_inst1.stoper_hc.measured_delay_hc_i_31\
        );

    \I__9987\ : InMux
    port map (
            O => \N__45768\,
            I => \N__45765\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__45765\,
            I => \N__45761\
        );

    \I__9985\ : InMux
    port map (
            O => \N__45764\,
            I => \N__45758\
        );

    \I__9984\ : Span4Mux_v
    port map (
            O => \N__45761\,
            I => \N__45753\
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__45758\,
            I => \N__45753\
        );

    \I__9982\ : Odrv4
    port map (
            O => \N__45753\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_1
        );

    \I__9981\ : InMux
    port map (
            O => \N__45750\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0\
        );

    \I__9980\ : InMux
    port map (
            O => \N__45747\,
            I => \N__45744\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__45744\,
            I => \N__45740\
        );

    \I__9978\ : InMux
    port map (
            O => \N__45743\,
            I => \N__45737\
        );

    \I__9977\ : Span4Mux_h
    port map (
            O => \N__45740\,
            I => \N__45734\
        );

    \I__9976\ : LocalMux
    port map (
            O => \N__45737\,
            I => \N__45731\
        );

    \I__9975\ : Odrv4
    port map (
            O => \N__45734\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_2
        );

    \I__9974\ : Odrv4
    port map (
            O => \N__45731\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_2
        );

    \I__9973\ : InMux
    port map (
            O => \N__45726\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1\
        );

    \I__9972\ : InMux
    port map (
            O => \N__45723\,
            I => \N__45719\
        );

    \I__9971\ : InMux
    port map (
            O => \N__45722\,
            I => \N__45716\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__45719\,
            I => \N__45713\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__45716\,
            I => \N__45710\
        );

    \I__9968\ : Odrv4
    port map (
            O => \N__45713\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_3
        );

    \I__9967\ : Odrv4
    port map (
            O => \N__45710\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_3
        );

    \I__9966\ : InMux
    port map (
            O => \N__45705\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2\
        );

    \I__9965\ : InMux
    port map (
            O => \N__45702\,
            I => \N__45698\
        );

    \I__9964\ : InMux
    port map (
            O => \N__45701\,
            I => \N__45695\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__45698\,
            I => \N__45692\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__45695\,
            I => \N__45689\
        );

    \I__9961\ : Odrv4
    port map (
            O => \N__45692\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_4
        );

    \I__9960\ : Odrv4
    port map (
            O => \N__45689\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_4
        );

    \I__9959\ : InMux
    port map (
            O => \N__45684\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3\
        );

    \I__9958\ : InMux
    port map (
            O => \N__45681\,
            I => \N__45678\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__45678\,
            I => \N__45675\
        );

    \I__9956\ : Span4Mux_s2_v
    port map (
            O => \N__45675\,
            I => \N__45672\
        );

    \I__9955\ : Span4Mux_v
    port map (
            O => \N__45672\,
            I => \N__45669\
        );

    \I__9954\ : Sp12to4
    port map (
            O => \N__45669\,
            I => \N__45666\
        );

    \I__9953\ : Span12Mux_h
    port map (
            O => \N__45666\,
            I => \N__45663\
        );

    \I__9952\ : Odrv12
    port map (
            O => \N__45663\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__9951\ : CascadeMux
    port map (
            O => \N__45660\,
            I => \N__45657\
        );

    \I__9950\ : InMux
    port map (
            O => \N__45657\,
            I => \N__45654\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__45654\,
            I => \N__45651\
        );

    \I__9948\ : Span4Mux_v
    port map (
            O => \N__45651\,
            I => \N__45648\
        );

    \I__9947\ : Sp12to4
    port map (
            O => \N__45648\,
            I => \N__45645\
        );

    \I__9946\ : Odrv12
    port map (
            O => \N__45645\,
            I => \pwm_generator_inst.un2_threshold_1_23\
        );

    \I__9945\ : InMux
    port map (
            O => \N__45642\,
            I => \N__45639\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__45639\,
            I => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\
        );

    \I__9943\ : InMux
    port map (
            O => \N__45636\,
            I => \bfn_16_29_0_\
        );

    \I__9942\ : InMux
    port map (
            O => \N__45633\,
            I => \N__45630\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__45630\,
            I => \N__45627\
        );

    \I__9940\ : Span4Mux_v
    port map (
            O => \N__45627\,
            I => \N__45624\
        );

    \I__9939\ : Span4Mux_h
    port map (
            O => \N__45624\,
            I => \N__45621\
        );

    \I__9938\ : Sp12to4
    port map (
            O => \N__45621\,
            I => \N__45618\
        );

    \I__9937\ : Span12Mux_h
    port map (
            O => \N__45618\,
            I => \N__45615\
        );

    \I__9936\ : Odrv12
    port map (
            O => \N__45615\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__9935\ : CascadeMux
    port map (
            O => \N__45612\,
            I => \N__45609\
        );

    \I__9934\ : InMux
    port map (
            O => \N__45609\,
            I => \N__45606\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__45606\,
            I => \N__45603\
        );

    \I__9932\ : Span4Mux_s3_v
    port map (
            O => \N__45603\,
            I => \N__45600\
        );

    \I__9931\ : Span4Mux_h
    port map (
            O => \N__45600\,
            I => \N__45597\
        );

    \I__9930\ : Span4Mux_h
    port map (
            O => \N__45597\,
            I => \N__45594\
        );

    \I__9929\ : Odrv4
    port map (
            O => \N__45594\,
            I => \pwm_generator_inst.un2_threshold_1_24\
        );

    \I__9928\ : InMux
    port map (
            O => \N__45591\,
            I => \N__45588\
        );

    \I__9927\ : LocalMux
    port map (
            O => \N__45588\,
            I => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\
        );

    \I__9926\ : InMux
    port map (
            O => \N__45585\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__9925\ : InMux
    port map (
            O => \N__45582\,
            I => \N__45579\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__45579\,
            I => \N__45576\
        );

    \I__9923\ : Span4Mux_s2_v
    port map (
            O => \N__45576\,
            I => \N__45573\
        );

    \I__9922\ : Span4Mux_v
    port map (
            O => \N__45573\,
            I => \N__45570\
        );

    \I__9921\ : Sp12to4
    port map (
            O => \N__45570\,
            I => \N__45567\
        );

    \I__9920\ : Span12Mux_h
    port map (
            O => \N__45567\,
            I => \N__45564\
        );

    \I__9919\ : Odrv12
    port map (
            O => \N__45564\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__9918\ : InMux
    port map (
            O => \N__45561\,
            I => \N__45558\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__45558\,
            I => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\
        );

    \I__9916\ : InMux
    port map (
            O => \N__45555\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__9915\ : CascadeMux
    port map (
            O => \N__45552\,
            I => \N__45549\
        );

    \I__9914\ : InMux
    port map (
            O => \N__45549\,
            I => \N__45546\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__45546\,
            I => \N__45543\
        );

    \I__9912\ : Sp12to4
    port map (
            O => \N__45543\,
            I => \N__45540\
        );

    \I__9911\ : Span12Mux_s6_v
    port map (
            O => \N__45540\,
            I => \N__45537\
        );

    \I__9910\ : Span12Mux_h
    port map (
            O => \N__45537\,
            I => \N__45534\
        );

    \I__9909\ : Odrv12
    port map (
            O => \N__45534\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__9908\ : InMux
    port map (
            O => \N__45531\,
            I => \N__45528\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__45528\,
            I => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\
        );

    \I__9906\ : InMux
    port map (
            O => \N__45525\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__9905\ : InMux
    port map (
            O => \N__45522\,
            I => \N__45519\
        );

    \I__9904\ : LocalMux
    port map (
            O => \N__45519\,
            I => \N__45516\
        );

    \I__9903\ : Span12Mux_s6_v
    port map (
            O => \N__45516\,
            I => \N__45513\
        );

    \I__9902\ : Span12Mux_h
    port map (
            O => \N__45513\,
            I => \N__45510\
        );

    \I__9901\ : Odrv12
    port map (
            O => \N__45510\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__9900\ : InMux
    port map (
            O => \N__45507\,
            I => \N__45504\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__45504\,
            I => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\
        );

    \I__9898\ : InMux
    port map (
            O => \N__45501\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__9897\ : CascadeMux
    port map (
            O => \N__45498\,
            I => \N__45495\
        );

    \I__9896\ : InMux
    port map (
            O => \N__45495\,
            I => \N__45492\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__45492\,
            I => \N__45489\
        );

    \I__9894\ : Span12Mux_h
    port map (
            O => \N__45489\,
            I => \N__45486\
        );

    \I__9893\ : Span12Mux_h
    port map (
            O => \N__45486\,
            I => \N__45483\
        );

    \I__9892\ : Odrv12
    port map (
            O => \N__45483\,
            I => \pwm_generator_inst.un2_threshold_2_13\
        );

    \I__9891\ : InMux
    port map (
            O => \N__45480\,
            I => \N__45477\
        );

    \I__9890\ : LocalMux
    port map (
            O => \N__45477\,
            I => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\
        );

    \I__9889\ : InMux
    port map (
            O => \N__45474\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12\
        );

    \I__9888\ : InMux
    port map (
            O => \N__45471\,
            I => \N__45468\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__45468\,
            I => \N__45465\
        );

    \I__9886\ : Span4Mux_s2_v
    port map (
            O => \N__45465\,
            I => \N__45462\
        );

    \I__9885\ : Span4Mux_v
    port map (
            O => \N__45462\,
            I => \N__45459\
        );

    \I__9884\ : Sp12to4
    port map (
            O => \N__45459\,
            I => \N__45456\
        );

    \I__9883\ : Span12Mux_h
    port map (
            O => \N__45456\,
            I => \N__45453\
        );

    \I__9882\ : Odrv12
    port map (
            O => \N__45453\,
            I => \pwm_generator_inst.un2_threshold_2_14\
        );

    \I__9881\ : InMux
    port map (
            O => \N__45450\,
            I => \N__45447\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__45447\,
            I => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\
        );

    \I__9879\ : InMux
    port map (
            O => \N__45444\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13\
        );

    \I__9878\ : InMux
    port map (
            O => \N__45441\,
            I => \N__45435\
        );

    \I__9877\ : CascadeMux
    port map (
            O => \N__45440\,
            I => \N__45431\
        );

    \I__9876\ : CascadeMux
    port map (
            O => \N__45439\,
            I => \N__45427\
        );

    \I__9875\ : CascadeMux
    port map (
            O => \N__45438\,
            I => \N__45423\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__45435\,
            I => \N__45420\
        );

    \I__9873\ : InMux
    port map (
            O => \N__45434\,
            I => \N__45407\
        );

    \I__9872\ : InMux
    port map (
            O => \N__45431\,
            I => \N__45407\
        );

    \I__9871\ : InMux
    port map (
            O => \N__45430\,
            I => \N__45407\
        );

    \I__9870\ : InMux
    port map (
            O => \N__45427\,
            I => \N__45407\
        );

    \I__9869\ : InMux
    port map (
            O => \N__45426\,
            I => \N__45407\
        );

    \I__9868\ : InMux
    port map (
            O => \N__45423\,
            I => \N__45407\
        );

    \I__9867\ : Span4Mux_v
    port map (
            O => \N__45420\,
            I => \N__45401\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__45407\,
            I => \N__45401\
        );

    \I__9865\ : InMux
    port map (
            O => \N__45406\,
            I => \N__45398\
        );

    \I__9864\ : Span4Mux_s2_v
    port map (
            O => \N__45401\,
            I => \N__45395\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__45398\,
            I => \N__45392\
        );

    \I__9862\ : Span4Mux_h
    port map (
            O => \N__45395\,
            I => \N__45389\
        );

    \I__9861\ : Span12Mux_h
    port map (
            O => \N__45392\,
            I => \N__45386\
        );

    \I__9860\ : Span4Mux_h
    port map (
            O => \N__45389\,
            I => \N__45383\
        );

    \I__9859\ : Odrv12
    port map (
            O => \N__45386\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__9858\ : Odrv4
    port map (
            O => \N__45383\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__9857\ : CascadeMux
    port map (
            O => \N__45378\,
            I => \N__45375\
        );

    \I__9856\ : InMux
    port map (
            O => \N__45375\,
            I => \N__45372\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__45372\,
            I => \N__45369\
        );

    \I__9854\ : Span4Mux_v
    port map (
            O => \N__45369\,
            I => \N__45366\
        );

    \I__9853\ : Odrv4
    port map (
            O => \N__45366\,
            I => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\
        );

    \I__9852\ : InMux
    port map (
            O => \N__45363\,
            I => \N__45360\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__45360\,
            I => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\
        );

    \I__9850\ : InMux
    port map (
            O => \N__45357\,
            I => \N__45354\
        );

    \I__9849\ : LocalMux
    port map (
            O => \N__45354\,
            I => \N__45351\
        );

    \I__9848\ : Span4Mux_h
    port map (
            O => \N__45351\,
            I => \N__45348\
        );

    \I__9847\ : Sp12to4
    port map (
            O => \N__45348\,
            I => \N__45345\
        );

    \I__9846\ : Span12Mux_s7_v
    port map (
            O => \N__45345\,
            I => \N__45342\
        );

    \I__9845\ : Span12Mux_h
    port map (
            O => \N__45342\,
            I => \N__45339\
        );

    \I__9844\ : Odrv12
    port map (
            O => \N__45339\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__9843\ : CascadeMux
    port map (
            O => \N__45336\,
            I => \N__45333\
        );

    \I__9842\ : InMux
    port map (
            O => \N__45333\,
            I => \N__45330\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__45330\,
            I => \N__45327\
        );

    \I__9840\ : Span4Mux_s3_v
    port map (
            O => \N__45327\,
            I => \N__45324\
        );

    \I__9839\ : Span4Mux_h
    port map (
            O => \N__45324\,
            I => \N__45321\
        );

    \I__9838\ : Span4Mux_h
    port map (
            O => \N__45321\,
            I => \N__45318\
        );

    \I__9837\ : Odrv4
    port map (
            O => \N__45318\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__9836\ : CascadeMux
    port map (
            O => \N__45315\,
            I => \N__45312\
        );

    \I__9835\ : InMux
    port map (
            O => \N__45312\,
            I => \N__45309\
        );

    \I__9834\ : LocalMux
    port map (
            O => \N__45309\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\
        );

    \I__9833\ : InMux
    port map (
            O => \N__45306\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__9832\ : InMux
    port map (
            O => \N__45303\,
            I => \N__45300\
        );

    \I__9831\ : LocalMux
    port map (
            O => \N__45300\,
            I => \N__45297\
        );

    \I__9830\ : Span4Mux_s3_v
    port map (
            O => \N__45297\,
            I => \N__45294\
        );

    \I__9829\ : Span4Mux_v
    port map (
            O => \N__45294\,
            I => \N__45291\
        );

    \I__9828\ : Sp12to4
    port map (
            O => \N__45291\,
            I => \N__45288\
        );

    \I__9827\ : Span12Mux_h
    port map (
            O => \N__45288\,
            I => \N__45285\
        );

    \I__9826\ : Odrv12
    port map (
            O => \N__45285\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__9825\ : CascadeMux
    port map (
            O => \N__45282\,
            I => \N__45279\
        );

    \I__9824\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45276\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__45276\,
            I => \N__45273\
        );

    \I__9822\ : Span4Mux_s3_v
    port map (
            O => \N__45273\,
            I => \N__45270\
        );

    \I__9821\ : Span4Mux_h
    port map (
            O => \N__45270\,
            I => \N__45267\
        );

    \I__9820\ : Span4Mux_h
    port map (
            O => \N__45267\,
            I => \N__45264\
        );

    \I__9819\ : Odrv4
    port map (
            O => \N__45264\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__9818\ : InMux
    port map (
            O => \N__45261\,
            I => \N__45258\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__45258\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\
        );

    \I__9816\ : InMux
    port map (
            O => \N__45255\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__9815\ : InMux
    port map (
            O => \N__45252\,
            I => \N__45249\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__45249\,
            I => \N__45246\
        );

    \I__9813\ : Span4Mux_h
    port map (
            O => \N__45246\,
            I => \N__45243\
        );

    \I__9812\ : Span4Mux_h
    port map (
            O => \N__45243\,
            I => \N__45240\
        );

    \I__9811\ : Span4Mux_h
    port map (
            O => \N__45240\,
            I => \N__45237\
        );

    \I__9810\ : Odrv4
    port map (
            O => \N__45237\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__9809\ : CascadeMux
    port map (
            O => \N__45234\,
            I => \N__45231\
        );

    \I__9808\ : InMux
    port map (
            O => \N__45231\,
            I => \N__45228\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__45228\,
            I => \N__45225\
        );

    \I__9806\ : Sp12to4
    port map (
            O => \N__45225\,
            I => \N__45222\
        );

    \I__9805\ : Span12Mux_s7_v
    port map (
            O => \N__45222\,
            I => \N__45219\
        );

    \I__9804\ : Span12Mux_h
    port map (
            O => \N__45219\,
            I => \N__45216\
        );

    \I__9803\ : Odrv12
    port map (
            O => \N__45216\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__9802\ : InMux
    port map (
            O => \N__45213\,
            I => \N__45210\
        );

    \I__9801\ : LocalMux
    port map (
            O => \N__45210\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\
        );

    \I__9800\ : InMux
    port map (
            O => \N__45207\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__9799\ : InMux
    port map (
            O => \N__45204\,
            I => \N__45201\
        );

    \I__9798\ : LocalMux
    port map (
            O => \N__45201\,
            I => \N__45198\
        );

    \I__9797\ : Span12Mux_s7_v
    port map (
            O => \N__45198\,
            I => \N__45195\
        );

    \I__9796\ : Span12Mux_h
    port map (
            O => \N__45195\,
            I => \N__45192\
        );

    \I__9795\ : Odrv12
    port map (
            O => \N__45192\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__9794\ : CascadeMux
    port map (
            O => \N__45189\,
            I => \N__45186\
        );

    \I__9793\ : InMux
    port map (
            O => \N__45186\,
            I => \N__45183\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__45183\,
            I => \N__45180\
        );

    \I__9791\ : Span12Mux_h
    port map (
            O => \N__45180\,
            I => \N__45177\
        );

    \I__9790\ : Odrv12
    port map (
            O => \N__45177\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__9789\ : InMux
    port map (
            O => \N__45174\,
            I => \N__45171\
        );

    \I__9788\ : LocalMux
    port map (
            O => \N__45171\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\
        );

    \I__9787\ : InMux
    port map (
            O => \N__45168\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__9786\ : InMux
    port map (
            O => \N__45165\,
            I => \N__45162\
        );

    \I__9785\ : LocalMux
    port map (
            O => \N__45162\,
            I => \N__45159\
        );

    \I__9784\ : Span12Mux_h
    port map (
            O => \N__45159\,
            I => \N__45156\
        );

    \I__9783\ : Span12Mux_h
    port map (
            O => \N__45156\,
            I => \N__45153\
        );

    \I__9782\ : Odrv12
    port map (
            O => \N__45153\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__9781\ : CascadeMux
    port map (
            O => \N__45150\,
            I => \N__45147\
        );

    \I__9780\ : InMux
    port map (
            O => \N__45147\,
            I => \N__45144\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__45144\,
            I => \N__45141\
        );

    \I__9778\ : Span4Mux_v
    port map (
            O => \N__45141\,
            I => \N__45138\
        );

    \I__9777\ : Sp12to4
    port map (
            O => \N__45138\,
            I => \N__45135\
        );

    \I__9776\ : Odrv12
    port map (
            O => \N__45135\,
            I => \pwm_generator_inst.un2_threshold_1_20\
        );

    \I__9775\ : InMux
    port map (
            O => \N__45132\,
            I => \N__45129\
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__45129\,
            I => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\
        );

    \I__9773\ : InMux
    port map (
            O => \N__45126\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__9772\ : InMux
    port map (
            O => \N__45123\,
            I => \N__45120\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__45120\,
            I => \N__45117\
        );

    \I__9770\ : Span4Mux_v
    port map (
            O => \N__45117\,
            I => \N__45114\
        );

    \I__9769\ : Span4Mux_h
    port map (
            O => \N__45114\,
            I => \N__45111\
        );

    \I__9768\ : Sp12to4
    port map (
            O => \N__45111\,
            I => \N__45108\
        );

    \I__9767\ : Span12Mux_h
    port map (
            O => \N__45108\,
            I => \N__45105\
        );

    \I__9766\ : Odrv12
    port map (
            O => \N__45105\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__9765\ : CascadeMux
    port map (
            O => \N__45102\,
            I => \N__45099\
        );

    \I__9764\ : InMux
    port map (
            O => \N__45099\,
            I => \N__45096\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__45096\,
            I => \N__45093\
        );

    \I__9762\ : Span12Mux_s5_v
    port map (
            O => \N__45093\,
            I => \N__45090\
        );

    \I__9761\ : Odrv12
    port map (
            O => \N__45090\,
            I => \pwm_generator_inst.un2_threshold_1_21\
        );

    \I__9760\ : InMux
    port map (
            O => \N__45087\,
            I => \N__45084\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__45084\,
            I => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\
        );

    \I__9758\ : InMux
    port map (
            O => \N__45081\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__9757\ : InMux
    port map (
            O => \N__45078\,
            I => \N__45075\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__45075\,
            I => \N__45072\
        );

    \I__9755\ : Span4Mux_h
    port map (
            O => \N__45072\,
            I => \N__45069\
        );

    \I__9754\ : Span4Mux_h
    port map (
            O => \N__45069\,
            I => \N__45066\
        );

    \I__9753\ : Sp12to4
    port map (
            O => \N__45066\,
            I => \N__45063\
        );

    \I__9752\ : Span12Mux_s7_v
    port map (
            O => \N__45063\,
            I => \N__45060\
        );

    \I__9751\ : Odrv12
    port map (
            O => \N__45060\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__9750\ : CascadeMux
    port map (
            O => \N__45057\,
            I => \N__45054\
        );

    \I__9749\ : InMux
    port map (
            O => \N__45054\,
            I => \N__45051\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__45051\,
            I => \N__45048\
        );

    \I__9747\ : Span4Mux_v
    port map (
            O => \N__45048\,
            I => \N__45045\
        );

    \I__9746\ : Sp12to4
    port map (
            O => \N__45045\,
            I => \N__45042\
        );

    \I__9745\ : Odrv12
    port map (
            O => \N__45042\,
            I => \pwm_generator_inst.un2_threshold_1_22\
        );

    \I__9744\ : InMux
    port map (
            O => \N__45039\,
            I => \N__45036\
        );

    \I__9743\ : LocalMux
    port map (
            O => \N__45036\,
            I => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\
        );

    \I__9742\ : InMux
    port map (
            O => \N__45033\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__9741\ : CascadeMux
    port map (
            O => \N__45030\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13_cascade_\
        );

    \I__9740\ : InMux
    port map (
            O => \N__45027\,
            I => \N__45023\
        );

    \I__9739\ : InMux
    port map (
            O => \N__45026\,
            I => \N__45020\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__45023\,
            I => \N__45015\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__45020\,
            I => \N__45015\
        );

    \I__9736\ : Odrv4
    port map (
            O => \N__45015\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__9735\ : InMux
    port map (
            O => \N__45012\,
            I => \N__45008\
        );

    \I__9734\ : InMux
    port map (
            O => \N__45011\,
            I => \N__45005\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__45008\,
            I => \N__45002\
        );

    \I__9732\ : LocalMux
    port map (
            O => \N__45005\,
            I => \N__44999\
        );

    \I__9731\ : Span4Mux_v
    port map (
            O => \N__45002\,
            I => \N__44996\
        );

    \I__9730\ : Span4Mux_v
    port map (
            O => \N__44999\,
            I => \N__44993\
        );

    \I__9729\ : Sp12to4
    port map (
            O => \N__44996\,
            I => \N__44990\
        );

    \I__9728\ : Span4Mux_h
    port map (
            O => \N__44993\,
            I => \N__44987\
        );

    \I__9727\ : Span12Mux_h
    port map (
            O => \N__44990\,
            I => \N__44982\
        );

    \I__9726\ : Sp12to4
    port map (
            O => \N__44987\,
            I => \N__44982\
        );

    \I__9725\ : Odrv12
    port map (
            O => \N__44982\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__9724\ : CascadeMux
    port map (
            O => \N__44979\,
            I => \N__44976\
        );

    \I__9723\ : InMux
    port map (
            O => \N__44976\,
            I => \N__44973\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__44973\,
            I => \N__44950\
        );

    \I__9721\ : InMux
    port map (
            O => \N__44972\,
            I => \N__44944\
        );

    \I__9720\ : InMux
    port map (
            O => \N__44971\,
            I => \N__44944\
        );

    \I__9719\ : InMux
    port map (
            O => \N__44970\,
            I => \N__44937\
        );

    \I__9718\ : InMux
    port map (
            O => \N__44969\,
            I => \N__44937\
        );

    \I__9717\ : InMux
    port map (
            O => \N__44968\,
            I => \N__44937\
        );

    \I__9716\ : InMux
    port map (
            O => \N__44967\,
            I => \N__44920\
        );

    \I__9715\ : InMux
    port map (
            O => \N__44966\,
            I => \N__44920\
        );

    \I__9714\ : InMux
    port map (
            O => \N__44965\,
            I => \N__44920\
        );

    \I__9713\ : InMux
    port map (
            O => \N__44964\,
            I => \N__44920\
        );

    \I__9712\ : InMux
    port map (
            O => \N__44963\,
            I => \N__44920\
        );

    \I__9711\ : InMux
    port map (
            O => \N__44962\,
            I => \N__44920\
        );

    \I__9710\ : InMux
    port map (
            O => \N__44961\,
            I => \N__44920\
        );

    \I__9709\ : InMux
    port map (
            O => \N__44960\,
            I => \N__44920\
        );

    \I__9708\ : InMux
    port map (
            O => \N__44959\,
            I => \N__44905\
        );

    \I__9707\ : InMux
    port map (
            O => \N__44958\,
            I => \N__44905\
        );

    \I__9706\ : InMux
    port map (
            O => \N__44957\,
            I => \N__44905\
        );

    \I__9705\ : InMux
    port map (
            O => \N__44956\,
            I => \N__44905\
        );

    \I__9704\ : InMux
    port map (
            O => \N__44955\,
            I => \N__44905\
        );

    \I__9703\ : InMux
    port map (
            O => \N__44954\,
            I => \N__44905\
        );

    \I__9702\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44905\
        );

    \I__9701\ : Span4Mux_v
    port map (
            O => \N__44950\,
            I => \N__44902\
        );

    \I__9700\ : InMux
    port map (
            O => \N__44949\,
            I => \N__44899\
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__44944\,
            I => \N__44894\
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__44937\,
            I => \N__44894\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__44920\,
            I => \N__44889\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__44905\,
            I => \N__44889\
        );

    \I__9695\ : Sp12to4
    port map (
            O => \N__44902\,
            I => \N__44882\
        );

    \I__9694\ : LocalMux
    port map (
            O => \N__44899\,
            I => \N__44882\
        );

    \I__9693\ : Span12Mux_s7_v
    port map (
            O => \N__44894\,
            I => \N__44882\
        );

    \I__9692\ : Span12Mux_s7_h
    port map (
            O => \N__44889\,
            I => \N__44879\
        );

    \I__9691\ : Span12Mux_h
    port map (
            O => \N__44882\,
            I => \N__44876\
        );

    \I__9690\ : Odrv12
    port map (
            O => \N__44879\,
            I => pwm_duty_input_10
        );

    \I__9689\ : Odrv12
    port map (
            O => \N__44876\,
            I => pwm_duty_input_10
        );

    \I__9688\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44868\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__44868\,
            I => \N__44865\
        );

    \I__9686\ : Span4Mux_v
    port map (
            O => \N__44865\,
            I => \N__44862\
        );

    \I__9685\ : Sp12to4
    port map (
            O => \N__44862\,
            I => \N__44859\
        );

    \I__9684\ : Span12Mux_h
    port map (
            O => \N__44859\,
            I => \N__44856\
        );

    \I__9683\ : Odrv12
    port map (
            O => \N__44856\,
            I => \pwm_generator_inst.un2_threshold_2_1_16\
        );

    \I__9682\ : InMux
    port map (
            O => \N__44853\,
            I => \N__44847\
        );

    \I__9681\ : InMux
    port map (
            O => \N__44852\,
            I => \N__44847\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__44847\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__9679\ : CascadeMux
    port map (
            O => \N__44844\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17_cascade_\
        );

    \I__9678\ : CascadeMux
    port map (
            O => \N__44841\,
            I => \N__44838\
        );

    \I__9677\ : InMux
    port map (
            O => \N__44838\,
            I => \N__44835\
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__44835\,
            I => \N__44831\
        );

    \I__9675\ : InMux
    port map (
            O => \N__44834\,
            I => \N__44828\
        );

    \I__9674\ : Odrv4
    port map (
            O => \N__44831\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__44828\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__9672\ : InMux
    port map (
            O => \N__44823\,
            I => \N__44820\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__44820\,
            I => \N__44817\
        );

    \I__9670\ : Span4Mux_s3_v
    port map (
            O => \N__44817\,
            I => \N__44814\
        );

    \I__9669\ : Span4Mux_v
    port map (
            O => \N__44814\,
            I => \N__44811\
        );

    \I__9668\ : Sp12to4
    port map (
            O => \N__44811\,
            I => \N__44808\
        );

    \I__9667\ : Span12Mux_h
    port map (
            O => \N__44808\,
            I => \N__44805\
        );

    \I__9666\ : Odrv12
    port map (
            O => \N__44805\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__9665\ : CascadeMux
    port map (
            O => \N__44802\,
            I => \N__44799\
        );

    \I__9664\ : InMux
    port map (
            O => \N__44799\,
            I => \N__44796\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__44796\,
            I => \N__44793\
        );

    \I__9662\ : Span4Mux_v
    port map (
            O => \N__44793\,
            I => \N__44790\
        );

    \I__9661\ : Sp12to4
    port map (
            O => \N__44790\,
            I => \N__44787\
        );

    \I__9660\ : Odrv12
    port map (
            O => \N__44787\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__9659\ : InMux
    port map (
            O => \N__44784\,
            I => \N__44781\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__44781\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_4\
        );

    \I__9657\ : InMux
    port map (
            O => \N__44778\,
            I => \bfn_16_24_0_\
        );

    \I__9656\ : InMux
    port map (
            O => \N__44775\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__9655\ : CascadeMux
    port map (
            O => \N__44772\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__9654\ : InMux
    port map (
            O => \N__44769\,
            I => \N__44766\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__44766\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__9652\ : CascadeMux
    port map (
            O => \N__44763\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__9651\ : InMux
    port map (
            O => \N__44760\,
            I => \N__44742\
        );

    \I__9650\ : InMux
    port map (
            O => \N__44759\,
            I => \N__44742\
        );

    \I__9649\ : InMux
    port map (
            O => \N__44758\,
            I => \N__44742\
        );

    \I__9648\ : InMux
    port map (
            O => \N__44757\,
            I => \N__44742\
        );

    \I__9647\ : InMux
    port map (
            O => \N__44756\,
            I => \N__44733\
        );

    \I__9646\ : InMux
    port map (
            O => \N__44755\,
            I => \N__44733\
        );

    \I__9645\ : InMux
    port map (
            O => \N__44754\,
            I => \N__44733\
        );

    \I__9644\ : InMux
    port map (
            O => \N__44753\,
            I => \N__44733\
        );

    \I__9643\ : InMux
    port map (
            O => \N__44752\,
            I => \N__44728\
        );

    \I__9642\ : InMux
    port map (
            O => \N__44751\,
            I => \N__44728\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__44742\,
            I => \N__44723\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__44733\,
            I => \N__44723\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__44728\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__9638\ : Odrv4
    port map (
            O => \N__44723\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__9637\ : CascadeMux
    port map (
            O => \N__44718\,
            I => \N__44715\
        );

    \I__9636\ : InMux
    port map (
            O => \N__44715\,
            I => \N__44712\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__44712\,
            I => \N__44708\
        );

    \I__9634\ : InMux
    port map (
            O => \N__44711\,
            I => \N__44705\
        );

    \I__9633\ : Odrv4
    port map (
            O => \N__44708\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__44705\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__9631\ : InMux
    port map (
            O => \N__44700\,
            I => \N__44694\
        );

    \I__9630\ : InMux
    port map (
            O => \N__44699\,
            I => \N__44694\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__44694\,
            I => \N__44691\
        );

    \I__9628\ : Odrv12
    port map (
            O => \N__44691\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__9627\ : InMux
    port map (
            O => \N__44688\,
            I => \N__44682\
        );

    \I__9626\ : InMux
    port map (
            O => \N__44687\,
            I => \N__44682\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__44682\,
            I => \N__44679\
        );

    \I__9624\ : Span4Mux_h
    port map (
            O => \N__44679\,
            I => \N__44676\
        );

    \I__9623\ : Odrv4
    port map (
            O => \N__44676\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__9622\ : CascadeMux
    port map (
            O => \N__44673\,
            I => \N__44670\
        );

    \I__9621\ : InMux
    port map (
            O => \N__44670\,
            I => \N__44664\
        );

    \I__9620\ : InMux
    port map (
            O => \N__44669\,
            I => \N__44664\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__44664\,
            I => \N__44661\
        );

    \I__9618\ : Span4Mux_h
    port map (
            O => \N__44661\,
            I => \N__44658\
        );

    \I__9617\ : Odrv4
    port map (
            O => \N__44658\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__9616\ : InMux
    port map (
            O => \N__44655\,
            I => \N__44652\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__44652\,
            I => \N__44649\
        );

    \I__9614\ : Span4Mux_v
    port map (
            O => \N__44649\,
            I => \N__44645\
        );

    \I__9613\ : InMux
    port map (
            O => \N__44648\,
            I => \N__44642\
        );

    \I__9612\ : Sp12to4
    port map (
            O => \N__44645\,
            I => \N__44637\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__44642\,
            I => \N__44637\
        );

    \I__9610\ : Odrv12
    port map (
            O => \N__44637\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__9609\ : InMux
    port map (
            O => \N__44634\,
            I => \N__44631\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__44631\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__9607\ : InMux
    port map (
            O => \N__44628\,
            I => \bfn_16_23_0_\
        );

    \I__9606\ : InMux
    port map (
            O => \N__44625\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__9605\ : InMux
    port map (
            O => \N__44622\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__9604\ : InMux
    port map (
            O => \N__44619\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__9603\ : InMux
    port map (
            O => \N__44616\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__9602\ : InMux
    port map (
            O => \N__44613\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__9601\ : InMux
    port map (
            O => \N__44610\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__9600\ : InMux
    port map (
            O => \N__44607\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__9599\ : CascadeMux
    port map (
            O => \N__44604\,
            I => \N__44600\
        );

    \I__9598\ : InMux
    port map (
            O => \N__44603\,
            I => \N__44597\
        );

    \I__9597\ : InMux
    port map (
            O => \N__44600\,
            I => \N__44594\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__44597\,
            I => \N__44591\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__44594\,
            I => \N__44588\
        );

    \I__9594\ : Span12Mux_s10_v
    port map (
            O => \N__44591\,
            I => \N__44585\
        );

    \I__9593\ : Span4Mux_h
    port map (
            O => \N__44588\,
            I => \N__44582\
        );

    \I__9592\ : Odrv12
    port map (
            O => \N__44585\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__9591\ : Odrv4
    port map (
            O => \N__44582\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__9590\ : InMux
    port map (
            O => \N__44577\,
            I => \N__44571\
        );

    \I__9589\ : InMux
    port map (
            O => \N__44576\,
            I => \N__44571\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__44571\,
            I => \N__44568\
        );

    \I__9587\ : Odrv12
    port map (
            O => \N__44568\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__9586\ : InMux
    port map (
            O => \N__44565\,
            I => \N__44559\
        );

    \I__9585\ : InMux
    port map (
            O => \N__44564\,
            I => \N__44559\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__44559\,
            I => \N__44556\
        );

    \I__9583\ : Odrv12
    port map (
            O => \N__44556\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__9582\ : InMux
    port map (
            O => \N__44553\,
            I => \N__44549\
        );

    \I__9581\ : InMux
    port map (
            O => \N__44552\,
            I => \N__44546\
        );

    \I__9580\ : LocalMux
    port map (
            O => \N__44549\,
            I => \N__44541\
        );

    \I__9579\ : LocalMux
    port map (
            O => \N__44546\,
            I => \N__44541\
        );

    \I__9578\ : Odrv12
    port map (
            O => \N__44541\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__9577\ : CascadeMux
    port map (
            O => \N__44538\,
            I => \N__44535\
        );

    \I__9576\ : InMux
    port map (
            O => \N__44535\,
            I => \N__44532\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__44532\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__9574\ : InMux
    port map (
            O => \N__44529\,
            I => \N__44523\
        );

    \I__9573\ : InMux
    port map (
            O => \N__44528\,
            I => \N__44523\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__44523\,
            I => \N__44520\
        );

    \I__9571\ : Span4Mux_h
    port map (
            O => \N__44520\,
            I => \N__44517\
        );

    \I__9570\ : Odrv4
    port map (
            O => \N__44517\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__9569\ : InMux
    port map (
            O => \N__44514\,
            I => \N__44511\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__44511\,
            I => \N__44507\
        );

    \I__9567\ : CascadeMux
    port map (
            O => \N__44510\,
            I => \N__44504\
        );

    \I__9566\ : Span4Mux_v
    port map (
            O => \N__44507\,
            I => \N__44501\
        );

    \I__9565\ : InMux
    port map (
            O => \N__44504\,
            I => \N__44498\
        );

    \I__9564\ : Sp12to4
    port map (
            O => \N__44501\,
            I => \N__44493\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__44498\,
            I => \N__44493\
        );

    \I__9562\ : Odrv12
    port map (
            O => \N__44493\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__9561\ : CascadeMux
    port map (
            O => \N__44490\,
            I => \N__44487\
        );

    \I__9560\ : InMux
    port map (
            O => \N__44487\,
            I => \N__44481\
        );

    \I__9559\ : InMux
    port map (
            O => \N__44486\,
            I => \N__44481\
        );

    \I__9558\ : LocalMux
    port map (
            O => \N__44481\,
            I => \N__44478\
        );

    \I__9557\ : Odrv12
    port map (
            O => \N__44478\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__9556\ : InMux
    port map (
            O => \N__44475\,
            I => \N__44472\
        );

    \I__9555\ : LocalMux
    port map (
            O => \N__44472\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\
        );

    \I__9554\ : InMux
    port map (
            O => \N__44469\,
            I => \N__44466\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__44466\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__9552\ : CascadeMux
    port map (
            O => \N__44463\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\
        );

    \I__9551\ : InMux
    port map (
            O => \N__44460\,
            I => \N__44457\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__44457\,
            I => \N__44454\
        );

    \I__9549\ : Span4Mux_v
    port map (
            O => \N__44454\,
            I => \N__44451\
        );

    \I__9548\ : Odrv4
    port map (
            O => \N__44451\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__9547\ : InMux
    port map (
            O => \N__44448\,
            I => \N__44445\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__44445\,
            I => \N__44441\
        );

    \I__9545\ : InMux
    port map (
            O => \N__44444\,
            I => \N__44438\
        );

    \I__9544\ : Span4Mux_h
    port map (
            O => \N__44441\,
            I => \N__44432\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__44438\,
            I => \N__44432\
        );

    \I__9542\ : InMux
    port map (
            O => \N__44437\,
            I => \N__44429\
        );

    \I__9541\ : Span4Mux_v
    port map (
            O => \N__44432\,
            I => \N__44425\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__44429\,
            I => \N__44422\
        );

    \I__9539\ : InMux
    port map (
            O => \N__44428\,
            I => \N__44419\
        );

    \I__9538\ : Sp12to4
    port map (
            O => \N__44425\,
            I => \N__44414\
        );

    \I__9537\ : Sp12to4
    port map (
            O => \N__44422\,
            I => \N__44414\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__44419\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__9535\ : Odrv12
    port map (
            O => \N__44414\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__9534\ : InMux
    port map (
            O => \N__44409\,
            I => \N__44406\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__44406\,
            I => \N__44403\
        );

    \I__9532\ : Span4Mux_v
    port map (
            O => \N__44403\,
            I => \N__44399\
        );

    \I__9531\ : InMux
    port map (
            O => \N__44402\,
            I => \N__44396\
        );

    \I__9530\ : Sp12to4
    port map (
            O => \N__44399\,
            I => \N__44391\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__44396\,
            I => \N__44391\
        );

    \I__9528\ : Odrv12
    port map (
            O => \N__44391\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__9527\ : CascadeMux
    port map (
            O => \N__44388\,
            I => \N__44384\
        );

    \I__9526\ : InMux
    port map (
            O => \N__44387\,
            I => \N__44381\
        );

    \I__9525\ : InMux
    port map (
            O => \N__44384\,
            I => \N__44378\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__44381\,
            I => \N__44375\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__44378\,
            I => \N__44372\
        );

    \I__9522\ : Span4Mux_h
    port map (
            O => \N__44375\,
            I => \N__44369\
        );

    \I__9521\ : Span12Mux_h
    port map (
            O => \N__44372\,
            I => \N__44366\
        );

    \I__9520\ : Span4Mux_h
    port map (
            O => \N__44369\,
            I => \N__44363\
        );

    \I__9519\ : Odrv12
    port map (
            O => \N__44366\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__9518\ : Odrv4
    port map (
            O => \N__44363\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__9517\ : CascadeMux
    port map (
            O => \N__44358\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\
        );

    \I__9516\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44352\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__44352\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__9514\ : InMux
    port map (
            O => \N__44349\,
            I => \N__44345\
        );

    \I__9513\ : InMux
    port map (
            O => \N__44348\,
            I => \N__44342\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__44345\,
            I => \N__44339\
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__44342\,
            I => \N__44336\
        );

    \I__9510\ : Span4Mux_h
    port map (
            O => \N__44339\,
            I => \N__44332\
        );

    \I__9509\ : Span4Mux_v
    port map (
            O => \N__44336\,
            I => \N__44329\
        );

    \I__9508\ : InMux
    port map (
            O => \N__44335\,
            I => \N__44326\
        );

    \I__9507\ : Span4Mux_h
    port map (
            O => \N__44332\,
            I => \N__44323\
        );

    \I__9506\ : Span4Mux_h
    port map (
            O => \N__44329\,
            I => \N__44320\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__44326\,
            I => \N__44317\
        );

    \I__9504\ : Span4Mux_h
    port map (
            O => \N__44323\,
            I => \N__44314\
        );

    \I__9503\ : Span4Mux_h
    port map (
            O => \N__44320\,
            I => \N__44311\
        );

    \I__9502\ : Span4Mux_h
    port map (
            O => \N__44317\,
            I => \N__44306\
        );

    \I__9501\ : Span4Mux_v
    port map (
            O => \N__44314\,
            I => \N__44306\
        );

    \I__9500\ : Odrv4
    port map (
            O => \N__44311\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__9499\ : Odrv4
    port map (
            O => \N__44306\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__9498\ : InMux
    port map (
            O => \N__44301\,
            I => \N__44298\
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__44298\,
            I => \N__44295\
        );

    \I__9496\ : Span4Mux_h
    port map (
            O => \N__44295\,
            I => \N__44292\
        );

    \I__9495\ : Span4Mux_v
    port map (
            O => \N__44292\,
            I => \N__44288\
        );

    \I__9494\ : InMux
    port map (
            O => \N__44291\,
            I => \N__44285\
        );

    \I__9493\ : Odrv4
    port map (
            O => \N__44288\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__44285\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__9491\ : InMux
    port map (
            O => \N__44280\,
            I => \N__44276\
        );

    \I__9490\ : InMux
    port map (
            O => \N__44279\,
            I => \N__44273\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__44276\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__44273\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__9487\ : InMux
    port map (
            O => \N__44268\,
            I => \N__44265\
        );

    \I__9486\ : LocalMux
    port map (
            O => \N__44265\,
            I => \N__44261\
        );

    \I__9485\ : InMux
    port map (
            O => \N__44264\,
            I => \N__44258\
        );

    \I__9484\ : Span4Mux_h
    port map (
            O => \N__44261\,
            I => \N__44255\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__44258\,
            I => \N__44252\
        );

    \I__9482\ : Span4Mux_v
    port map (
            O => \N__44255\,
            I => \N__44249\
        );

    \I__9481\ : Span4Mux_v
    port map (
            O => \N__44252\,
            I => \N__44246\
        );

    \I__9480\ : Odrv4
    port map (
            O => \N__44249\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__9479\ : Odrv4
    port map (
            O => \N__44246\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__9478\ : InMux
    port map (
            O => \N__44241\,
            I => \N__44237\
        );

    \I__9477\ : InMux
    port map (
            O => \N__44240\,
            I => \N__44234\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__44237\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__44234\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__9474\ : InMux
    port map (
            O => \N__44229\,
            I => \N__44225\
        );

    \I__9473\ : InMux
    port map (
            O => \N__44228\,
            I => \N__44222\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__44225\,
            I => \N__44219\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__44222\,
            I => \N__44216\
        );

    \I__9470\ : Span4Mux_v
    port map (
            O => \N__44219\,
            I => \N__44213\
        );

    \I__9469\ : Span4Mux_v
    port map (
            O => \N__44216\,
            I => \N__44208\
        );

    \I__9468\ : Span4Mux_h
    port map (
            O => \N__44213\,
            I => \N__44208\
        );

    \I__9467\ : Odrv4
    port map (
            O => \N__44208\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__9466\ : CascadeMux
    port map (
            O => \N__44205\,
            I => \N__44202\
        );

    \I__9465\ : InMux
    port map (
            O => \N__44202\,
            I => \N__44198\
        );

    \I__9464\ : InMux
    port map (
            O => \N__44201\,
            I => \N__44195\
        );

    \I__9463\ : LocalMux
    port map (
            O => \N__44198\,
            I => \N__44192\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__44195\,
            I => \N__44189\
        );

    \I__9461\ : Span4Mux_v
    port map (
            O => \N__44192\,
            I => \N__44184\
        );

    \I__9460\ : Span4Mux_h
    port map (
            O => \N__44189\,
            I => \N__44184\
        );

    \I__9459\ : Odrv4
    port map (
            O => \N__44184\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__9458\ : CascadeMux
    port map (
            O => \N__44181\,
            I => \N__44178\
        );

    \I__9457\ : InMux
    port map (
            O => \N__44178\,
            I => \N__44174\
        );

    \I__9456\ : InMux
    port map (
            O => \N__44177\,
            I => \N__44171\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__44174\,
            I => \N__44168\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__44171\,
            I => \N__44165\
        );

    \I__9453\ : Span4Mux_v
    port map (
            O => \N__44168\,
            I => \N__44162\
        );

    \I__9452\ : Span4Mux_v
    port map (
            O => \N__44165\,
            I => \N__44157\
        );

    \I__9451\ : Span4Mux_h
    port map (
            O => \N__44162\,
            I => \N__44157\
        );

    \I__9450\ : Odrv4
    port map (
            O => \N__44157\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__9449\ : InMux
    port map (
            O => \N__44154\,
            I => \N__44150\
        );

    \I__9448\ : InMux
    port map (
            O => \N__44153\,
            I => \N__44147\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__44150\,
            I => \N__44144\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__44147\,
            I => \N__44141\
        );

    \I__9445\ : Span4Mux_h
    port map (
            O => \N__44144\,
            I => \N__44138\
        );

    \I__9444\ : Odrv12
    port map (
            O => \N__44141\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__9443\ : Odrv4
    port map (
            O => \N__44138\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__9442\ : InMux
    port map (
            O => \N__44133\,
            I => \N__44130\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__44130\,
            I => \N__44127\
        );

    \I__9440\ : Span4Mux_h
    port map (
            O => \N__44127\,
            I => \N__44124\
        );

    \I__9439\ : Span4Mux_v
    port map (
            O => \N__44124\,
            I => \N__44120\
        );

    \I__9438\ : InMux
    port map (
            O => \N__44123\,
            I => \N__44117\
        );

    \I__9437\ : Odrv4
    port map (
            O => \N__44120\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__44117\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__9435\ : InMux
    port map (
            O => \N__44112\,
            I => \N__44087\
        );

    \I__9434\ : InMux
    port map (
            O => \N__44111\,
            I => \N__44087\
        );

    \I__9433\ : InMux
    port map (
            O => \N__44110\,
            I => \N__44078\
        );

    \I__9432\ : InMux
    port map (
            O => \N__44109\,
            I => \N__44078\
        );

    \I__9431\ : InMux
    port map (
            O => \N__44108\,
            I => \N__44078\
        );

    \I__9430\ : InMux
    port map (
            O => \N__44107\,
            I => \N__44078\
        );

    \I__9429\ : InMux
    port map (
            O => \N__44106\,
            I => \N__44075\
        );

    \I__9428\ : InMux
    port map (
            O => \N__44105\,
            I => \N__44066\
        );

    \I__9427\ : InMux
    port map (
            O => \N__44104\,
            I => \N__44061\
        );

    \I__9426\ : InMux
    port map (
            O => \N__44103\,
            I => \N__44061\
        );

    \I__9425\ : InMux
    port map (
            O => \N__44102\,
            I => \N__44054\
        );

    \I__9424\ : InMux
    port map (
            O => \N__44101\,
            I => \N__44054\
        );

    \I__9423\ : InMux
    port map (
            O => \N__44100\,
            I => \N__44054\
        );

    \I__9422\ : InMux
    port map (
            O => \N__44099\,
            I => \N__44051\
        );

    \I__9421\ : InMux
    port map (
            O => \N__44098\,
            I => \N__44048\
        );

    \I__9420\ : InMux
    port map (
            O => \N__44097\,
            I => \N__44045\
        );

    \I__9419\ : InMux
    port map (
            O => \N__44096\,
            I => \N__44037\
        );

    \I__9418\ : InMux
    port map (
            O => \N__44095\,
            I => \N__44037\
        );

    \I__9417\ : InMux
    port map (
            O => \N__44094\,
            I => \N__44030\
        );

    \I__9416\ : InMux
    port map (
            O => \N__44093\,
            I => \N__44030\
        );

    \I__9415\ : InMux
    port map (
            O => \N__44092\,
            I => \N__44030\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__44087\,
            I => \N__44023\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__44078\,
            I => \N__44023\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__44075\,
            I => \N__44023\
        );

    \I__9411\ : InMux
    port map (
            O => \N__44074\,
            I => \N__44020\
        );

    \I__9410\ : InMux
    port map (
            O => \N__44073\,
            I => \N__44009\
        );

    \I__9409\ : InMux
    port map (
            O => \N__44072\,
            I => \N__44009\
        );

    \I__9408\ : InMux
    port map (
            O => \N__44071\,
            I => \N__44009\
        );

    \I__9407\ : InMux
    port map (
            O => \N__44070\,
            I => \N__44009\
        );

    \I__9406\ : InMux
    port map (
            O => \N__44069\,
            I => \N__44009\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__44066\,
            I => \N__44002\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__44061\,
            I => \N__44002\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__44054\,
            I => \N__44002\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__44051\,
            I => \N__43995\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__44048\,
            I => \N__43995\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__44045\,
            I => \N__43995\
        );

    \I__9399\ : InMux
    port map (
            O => \N__44044\,
            I => \N__43990\
        );

    \I__9398\ : InMux
    port map (
            O => \N__44043\,
            I => \N__43990\
        );

    \I__9397\ : InMux
    port map (
            O => \N__44042\,
            I => \N__43987\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__44037\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__44030\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__9394\ : Odrv12
    port map (
            O => \N__44023\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__44020\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__44009\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__9391\ : Odrv4
    port map (
            O => \N__44002\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__9390\ : Odrv4
    port map (
            O => \N__43995\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__43990\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__43987\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__9387\ : InMux
    port map (
            O => \N__43968\,
            I => \N__43964\
        );

    \I__9386\ : InMux
    port map (
            O => \N__43967\,
            I => \N__43961\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__43964\,
            I => \N__43958\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__43961\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__9383\ : Odrv4
    port map (
            O => \N__43958\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__9382\ : InMux
    port map (
            O => \N__43953\,
            I => \N__43949\
        );

    \I__9381\ : InMux
    port map (
            O => \N__43952\,
            I => \N__43946\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__43949\,
            I => \N__43943\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__43946\,
            I => \N__43940\
        );

    \I__9378\ : Span4Mux_h
    port map (
            O => \N__43943\,
            I => \N__43937\
        );

    \I__9377\ : Odrv12
    port map (
            O => \N__43940\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__9376\ : Odrv4
    port map (
            O => \N__43937\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__9375\ : InMux
    port map (
            O => \N__43932\,
            I => \N__43928\
        );

    \I__9374\ : InMux
    port map (
            O => \N__43931\,
            I => \N__43925\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__43928\,
            I => \N__43922\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__43925\,
            I => \N__43919\
        );

    \I__9371\ : Span4Mux_h
    port map (
            O => \N__43922\,
            I => \N__43916\
        );

    \I__9370\ : Odrv12
    port map (
            O => \N__43919\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__9369\ : Odrv4
    port map (
            O => \N__43916\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__9368\ : InMux
    port map (
            O => \N__43911\,
            I => \N__43908\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__43908\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__9366\ : InMux
    port map (
            O => \N__43905\,
            I => \N__43902\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__43902\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__9364\ : InMux
    port map (
            O => \N__43899\,
            I => \N__43896\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__43896\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__9362\ : CascadeMux
    port map (
            O => \N__43893\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\
        );

    \I__9361\ : InMux
    port map (
            O => \N__43890\,
            I => \N__43887\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__43887\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\
        );

    \I__9359\ : CascadeMux
    port map (
            O => \N__43884\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_\
        );

    \I__9358\ : CascadeMux
    port map (
            O => \N__43881\,
            I => \N__43878\
        );

    \I__9357\ : InMux
    port map (
            O => \N__43878\,
            I => \N__43875\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__43875\,
            I => \N__43872\
        );

    \I__9355\ : Odrv4
    port map (
            O => \N__43872\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\
        );

    \I__9354\ : InMux
    port map (
            O => \N__43869\,
            I => \N__43866\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__43866\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\
        );

    \I__9352\ : InMux
    port map (
            O => \N__43863\,
            I => \N__43859\
        );

    \I__9351\ : CascadeMux
    port map (
            O => \N__43862\,
            I => \N__43856\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__43859\,
            I => \N__43853\
        );

    \I__9349\ : InMux
    port map (
            O => \N__43856\,
            I => \N__43850\
        );

    \I__9348\ : Span4Mux_h
    port map (
            O => \N__43853\,
            I => \N__43845\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__43850\,
            I => \N__43845\
        );

    \I__9346\ : Span4Mux_v
    port map (
            O => \N__43845\,
            I => \N__43842\
        );

    \I__9345\ : Odrv4
    port map (
            O => \N__43842\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__9344\ : InMux
    port map (
            O => \N__43839\,
            I => \N__43836\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__43836\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__9342\ : CascadeMux
    port map (
            O => \N__43833\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4_cascade_\
        );

    \I__9341\ : InMux
    port map (
            O => \N__43830\,
            I => \N__43827\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__43827\,
            I => \N__43824\
        );

    \I__9339\ : Span4Mux_v
    port map (
            O => \N__43824\,
            I => \N__43821\
        );

    \I__9338\ : Odrv4
    port map (
            O => \N__43821\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4\
        );

    \I__9337\ : InMux
    port map (
            O => \N__43818\,
            I => \N__43815\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__43815\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\
        );

    \I__9335\ : InMux
    port map (
            O => \N__43812\,
            I => \N__43808\
        );

    \I__9334\ : InMux
    port map (
            O => \N__43811\,
            I => \N__43805\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__43808\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__43805\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__9331\ : InMux
    port map (
            O => \N__43800\,
            I => \N__43796\
        );

    \I__9330\ : InMux
    port map (
            O => \N__43799\,
            I => \N__43793\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__43796\,
            I => \N__43790\
        );

    \I__9328\ : LocalMux
    port map (
            O => \N__43793\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__9327\ : Odrv4
    port map (
            O => \N__43790\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__9326\ : InMux
    port map (
            O => \N__43785\,
            I => \N__43781\
        );

    \I__9325\ : InMux
    port map (
            O => \N__43784\,
            I => \N__43778\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__43781\,
            I => \N__43775\
        );

    \I__9323\ : LocalMux
    port map (
            O => \N__43778\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__9322\ : Odrv12
    port map (
            O => \N__43775\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__9321\ : InMux
    port map (
            O => \N__43770\,
            I => \N__43767\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__43767\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__9319\ : CascadeMux
    port map (
            O => \N__43764\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\
        );

    \I__9318\ : CascadeMux
    port map (
            O => \N__43761\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\
        );

    \I__9317\ : InMux
    port map (
            O => \N__43758\,
            I => \N__43755\
        );

    \I__9316\ : LocalMux
    port map (
            O => \N__43755\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\
        );

    \I__9315\ : InMux
    port map (
            O => \N__43752\,
            I => \N__43749\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__43749\,
            I => \N__43746\
        );

    \I__9313\ : Span4Mux_h
    port map (
            O => \N__43746\,
            I => \N__43742\
        );

    \I__9312\ : CascadeMux
    port map (
            O => \N__43745\,
            I => \N__43739\
        );

    \I__9311\ : Span4Mux_v
    port map (
            O => \N__43742\,
            I => \N__43736\
        );

    \I__9310\ : InMux
    port map (
            O => \N__43739\,
            I => \N__43733\
        );

    \I__9309\ : Odrv4
    port map (
            O => \N__43736\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__43733\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9307\ : InMux
    port map (
            O => \N__43728\,
            I => \N__43725\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__43725\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__9305\ : CascadeMux
    port map (
            O => \N__43722\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\
        );

    \I__9304\ : InMux
    port map (
            O => \N__43719\,
            I => \N__43716\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__43716\,
            I => \N__43713\
        );

    \I__9302\ : Span4Mux_v
    port map (
            O => \N__43713\,
            I => \N__43710\
        );

    \I__9301\ : Odrv4
    port map (
            O => \N__43710\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15\
        );

    \I__9300\ : CascadeMux
    port map (
            O => \N__43707\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\
        );

    \I__9299\ : InMux
    port map (
            O => \N__43704\,
            I => \N__43698\
        );

    \I__9298\ : InMux
    port map (
            O => \N__43703\,
            I => \N__43698\
        );

    \I__9297\ : LocalMux
    port map (
            O => \N__43698\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__9296\ : InMux
    port map (
            O => \N__43695\,
            I => \N__43692\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__43692\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__9294\ : CascadeMux
    port map (
            O => \N__43689\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11_cascade_\
        );

    \I__9293\ : InMux
    port map (
            O => \N__43686\,
            I => \N__43683\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__43683\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__9291\ : CascadeMux
    port map (
            O => \N__43680\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\
        );

    \I__9290\ : CascadeMux
    port map (
            O => \N__43677\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\
        );

    \I__9289\ : InMux
    port map (
            O => \N__43674\,
            I => \N__43670\
        );

    \I__9288\ : InMux
    port map (
            O => \N__43673\,
            I => \N__43667\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__43670\,
            I => \N__43664\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__43667\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__9285\ : Odrv12
    port map (
            O => \N__43664\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__9284\ : InMux
    port map (
            O => \N__43659\,
            I => \N__43655\
        );

    \I__9283\ : InMux
    port map (
            O => \N__43658\,
            I => \N__43652\
        );

    \I__9282\ : LocalMux
    port map (
            O => \N__43655\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__43652\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__9280\ : CascadeMux
    port map (
            O => \N__43647\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16_cascade_\
        );

    \I__9279\ : InMux
    port map (
            O => \N__43644\,
            I => \N__43641\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__43641\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__9277\ : CascadeMux
    port map (
            O => \N__43638\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\
        );

    \I__9276\ : InMux
    port map (
            O => \N__43635\,
            I => \N__43632\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__43632\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__9274\ : CascadeMux
    port map (
            O => \N__43629\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4_cascade_\
        );

    \I__9273\ : InMux
    port map (
            O => \N__43626\,
            I => \N__43623\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__43623\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__9271\ : CascadeMux
    port map (
            O => \N__43620\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15_cascade_\
        );

    \I__9270\ : InMux
    port map (
            O => \N__43617\,
            I => \N__43614\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__43614\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__9268\ : InMux
    port map (
            O => \N__43611\,
            I => \N__43608\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__43608\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__9266\ : CascadeMux
    port map (
            O => \N__43605\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\
        );

    \I__9265\ : InMux
    port map (
            O => \N__43602\,
            I => \N__43599\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__43599\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__9263\ : CascadeMux
    port map (
            O => \N__43596\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3_cascade_\
        );

    \I__9262\ : InMux
    port map (
            O => \N__43593\,
            I => \N__43590\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__43590\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__9260\ : CascadeMux
    port map (
            O => \N__43587\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\
        );

    \I__9259\ : InMux
    port map (
            O => \N__43584\,
            I => \N__43581\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__43581\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__9257\ : CascadeMux
    port map (
            O => \N__43578\,
            I => \N__43575\
        );

    \I__9256\ : InMux
    port map (
            O => \N__43575\,
            I => \N__43569\
        );

    \I__9255\ : InMux
    port map (
            O => \N__43574\,
            I => \N__43569\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__43569\,
            I => \N__43566\
        );

    \I__9253\ : Span4Mux_v
    port map (
            O => \N__43566\,
            I => \N__43563\
        );

    \I__9252\ : Odrv4
    port map (
            O => \N__43563\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_26\
        );

    \I__9251\ : InMux
    port map (
            O => \N__43560\,
            I => \N__43554\
        );

    \I__9250\ : InMux
    port map (
            O => \N__43559\,
            I => \N__43554\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__43554\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_21\
        );

    \I__9248\ : InMux
    port map (
            O => \N__43551\,
            I => \N__43548\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__43548\,
            I => \N__43545\
        );

    \I__9246\ : Span4Mux_h
    port map (
            O => \N__43545\,
            I => \N__43542\
        );

    \I__9245\ : Odrv4
    port map (
            O => \N__43542\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_4\
        );

    \I__9244\ : InMux
    port map (
            O => \N__43539\,
            I => \N__43533\
        );

    \I__9243\ : InMux
    port map (
            O => \N__43538\,
            I => \N__43533\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__43533\,
            I => \N__43530\
        );

    \I__9241\ : Odrv4
    port map (
            O => \N__43530\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_16\
        );

    \I__9240\ : InMux
    port map (
            O => \N__43527\,
            I => \N__43521\
        );

    \I__9239\ : InMux
    port map (
            O => \N__43526\,
            I => \N__43521\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__43521\,
            I => \N__43518\
        );

    \I__9237\ : Odrv4
    port map (
            O => \N__43518\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_19\
        );

    \I__9236\ : InMux
    port map (
            O => \N__43515\,
            I => \N__43512\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__43512\,
            I => \N__43509\
        );

    \I__9234\ : Span4Mux_v
    port map (
            O => \N__43509\,
            I => \N__43506\
        );

    \I__9233\ : Sp12to4
    port map (
            O => \N__43506\,
            I => \N__43503\
        );

    \I__9232\ : Odrv12
    port map (
            O => \N__43503\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_7\
        );

    \I__9231\ : InMux
    port map (
            O => \N__43500\,
            I => \N__43496\
        );

    \I__9230\ : InMux
    port map (
            O => \N__43499\,
            I => \N__43493\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__43496\,
            I => \N__43490\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__43493\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24\
        );

    \I__9227\ : Odrv4
    port map (
            O => \N__43490\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24\
        );

    \I__9226\ : InMux
    port map (
            O => \N__43485\,
            I => \N__43481\
        );

    \I__9225\ : InMux
    port map (
            O => \N__43484\,
            I => \N__43478\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__43481\,
            I => \N__43475\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__43478\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25\
        );

    \I__9222\ : Odrv4
    port map (
            O => \N__43475\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25\
        );

    \I__9221\ : CEMux
    port map (
            O => \N__43470\,
            I => \N__43463\
        );

    \I__9220\ : CEMux
    port map (
            O => \N__43469\,
            I => \N__43460\
        );

    \I__9219\ : CEMux
    port map (
            O => \N__43468\,
            I => \N__43457\
        );

    \I__9218\ : CEMux
    port map (
            O => \N__43467\,
            I => \N__43453\
        );

    \I__9217\ : CEMux
    port map (
            O => \N__43466\,
            I => \N__43450\
        );

    \I__9216\ : LocalMux
    port map (
            O => \N__43463\,
            I => \N__43445\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__43460\,
            I => \N__43445\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__43457\,
            I => \N__43442\
        );

    \I__9213\ : CEMux
    port map (
            O => \N__43456\,
            I => \N__43439\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__43453\,
            I => \N__43436\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__43450\,
            I => \N__43432\
        );

    \I__9210\ : Span4Mux_v
    port map (
            O => \N__43445\,
            I => \N__43425\
        );

    \I__9209\ : Span4Mux_v
    port map (
            O => \N__43442\,
            I => \N__43425\
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__43439\,
            I => \N__43425\
        );

    \I__9207\ : Span4Mux_v
    port map (
            O => \N__43436\,
            I => \N__43422\
        );

    \I__9206\ : CEMux
    port map (
            O => \N__43435\,
            I => \N__43419\
        );

    \I__9205\ : Span4Mux_v
    port map (
            O => \N__43432\,
            I => \N__43416\
        );

    \I__9204\ : Span4Mux_v
    port map (
            O => \N__43425\,
            I => \N__43413\
        );

    \I__9203\ : Span4Mux_v
    port map (
            O => \N__43422\,
            I => \N__43408\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__43419\,
            I => \N__43408\
        );

    \I__9201\ : Span4Mux_v
    port map (
            O => \N__43416\,
            I => \N__43405\
        );

    \I__9200\ : Span4Mux_h
    port map (
            O => \N__43413\,
            I => \N__43402\
        );

    \I__9199\ : Span4Mux_h
    port map (
            O => \N__43408\,
            I => \N__43399\
        );

    \I__9198\ : Odrv4
    port map (
            O => \N__43405\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__9197\ : Odrv4
    port map (
            O => \N__43402\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__9196\ : Odrv4
    port map (
            O => \N__43399\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__9195\ : InMux
    port map (
            O => \N__43392\,
            I => \N__43389\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__43389\,
            I => \N__43386\
        );

    \I__9193\ : Odrv4
    port map (
            O => \N__43386\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_13\
        );

    \I__9192\ : InMux
    port map (
            O => \N__43383\,
            I => \N__43380\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__43380\,
            I => \N__43377\
        );

    \I__9190\ : Odrv4
    port map (
            O => \N__43377\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_8\
        );

    \I__9189\ : InMux
    port map (
            O => \N__43374\,
            I => \N__43371\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__43371\,
            I => \N__43368\
        );

    \I__9187\ : Span4Mux_h
    port map (
            O => \N__43368\,
            I => \N__43365\
        );

    \I__9186\ : Odrv4
    port map (
            O => \N__43365\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_3\
        );

    \I__9185\ : InMux
    port map (
            O => \N__43362\,
            I => \N__43359\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__43359\,
            I => \N__43356\
        );

    \I__9183\ : Span4Mux_v
    port map (
            O => \N__43356\,
            I => \N__43353\
        );

    \I__9182\ : Odrv4
    port map (
            O => \N__43353\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_15\
        );

    \I__9181\ : InMux
    port map (
            O => \N__43350\,
            I => \N__43347\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__43347\,
            I => \N__43344\
        );

    \I__9179\ : Span4Mux_v
    port map (
            O => \N__43344\,
            I => \N__43341\
        );

    \I__9178\ : Odrv4
    port map (
            O => \N__43341\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_5\
        );

    \I__9177\ : InMux
    port map (
            O => \N__43338\,
            I => \N__43335\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__43335\,
            I => \N__43332\
        );

    \I__9175\ : Span4Mux_h
    port map (
            O => \N__43332\,
            I => \N__43329\
        );

    \I__9174\ : Odrv4
    port map (
            O => \N__43329\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_13\
        );

    \I__9173\ : InMux
    port map (
            O => \N__43326\,
            I => \N__43323\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__43323\,
            I => \N__43320\
        );

    \I__9171\ : Span4Mux_h
    port map (
            O => \N__43320\,
            I => \N__43317\
        );

    \I__9170\ : Odrv4
    port map (
            O => \N__43317\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_14\
        );

    \I__9169\ : CascadeMux
    port map (
            O => \N__43314\,
            I => \N__43310\
        );

    \I__9168\ : InMux
    port map (
            O => \N__43313\,
            I => \N__43305\
        );

    \I__9167\ : InMux
    port map (
            O => \N__43310\,
            I => \N__43305\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__43305\,
            I => \N__43302\
        );

    \I__9165\ : Span12Mux_h
    port map (
            O => \N__43302\,
            I => \N__43299\
        );

    \I__9164\ : Odrv12
    port map (
            O => \N__43299\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_27\
        );

    \I__9163\ : InMux
    port map (
            O => \N__43296\,
            I => \N__43293\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__43293\,
            I => \N__43290\
        );

    \I__9161\ : Span4Mux_h
    port map (
            O => \N__43290\,
            I => \N__43287\
        );

    \I__9160\ : Odrv4
    port map (
            O => \N__43287\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_9\
        );

    \I__9159\ : InMux
    port map (
            O => \N__43284\,
            I => \N__43281\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__43281\,
            I => \N__43278\
        );

    \I__9157\ : Span4Mux_h
    port map (
            O => \N__43278\,
            I => \N__43275\
        );

    \I__9156\ : Odrv4
    port map (
            O => \N__43275\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_10\
        );

    \I__9155\ : InMux
    port map (
            O => \N__43272\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__9154\ : InMux
    port map (
            O => \N__43269\,
            I => \N__43266\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__43266\,
            I => \N__43263\
        );

    \I__9152\ : Span4Mux_h
    port map (
            O => \N__43263\,
            I => \N__43260\
        );

    \I__9151\ : Odrv4
    port map (
            O => \N__43260\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_11\
        );

    \I__9150\ : InMux
    port map (
            O => \N__43257\,
            I => \N__43254\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__43254\,
            I => \N__43251\
        );

    \I__9148\ : Span4Mux_h
    port map (
            O => \N__43251\,
            I => \N__43248\
        );

    \I__9147\ : Odrv4
    port map (
            O => \N__43248\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_14\
        );

    \I__9146\ : InMux
    port map (
            O => \N__43245\,
            I => \N__43242\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__43242\,
            I => \N__43239\
        );

    \I__9144\ : Odrv4
    port map (
            O => \N__43239\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_5\
        );

    \I__9143\ : InMux
    port map (
            O => \N__43236\,
            I => \N__43233\
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__43233\,
            I => \N__43230\
        );

    \I__9141\ : Odrv4
    port map (
            O => \N__43230\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_7\
        );

    \I__9140\ : InMux
    port map (
            O => \N__43227\,
            I => \N__43224\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__43224\,
            I => \N__43221\
        );

    \I__9138\ : Odrv4
    port map (
            O => \N__43221\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_10\
        );

    \I__9137\ : InMux
    port map (
            O => \N__43218\,
            I => \N__43215\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__43215\,
            I => \N__43212\
        );

    \I__9135\ : Odrv4
    port map (
            O => \N__43212\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_15\
        );

    \I__9134\ : InMux
    port map (
            O => \N__43209\,
            I => \N__43206\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__43206\,
            I => \N__43203\
        );

    \I__9132\ : Odrv4
    port map (
            O => \N__43203\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_12\
        );

    \I__9131\ : InMux
    port map (
            O => \N__43200\,
            I => \N__43197\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__43197\,
            I => \N__43194\
        );

    \I__9129\ : Odrv4
    port map (
            O => \N__43194\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_9\
        );

    \I__9128\ : InMux
    port map (
            O => \N__43191\,
            I => \N__43188\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__43188\,
            I => \N__43185\
        );

    \I__9126\ : Span4Mux_v
    port map (
            O => \N__43185\,
            I => \N__43182\
        );

    \I__9125\ : Sp12to4
    port map (
            O => \N__43182\,
            I => \N__43179\
        );

    \I__9124\ : Odrv12
    port map (
            O => \N__43179\,
            I => \pwm_generator_inst.O_13\
        );

    \I__9123\ : InMux
    port map (
            O => \N__43176\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__9122\ : InMux
    port map (
            O => \N__43173\,
            I => \N__43170\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__43170\,
            I => \N__43167\
        );

    \I__9120\ : Span12Mux_s6_v
    port map (
            O => \N__43167\,
            I => \N__43164\
        );

    \I__9119\ : Odrv12
    port map (
            O => \N__43164\,
            I => \pwm_generator_inst.O_14\
        );

    \I__9118\ : InMux
    port map (
            O => \N__43161\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__9117\ : InMux
    port map (
            O => \N__43158\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__9116\ : InMux
    port map (
            O => \N__43155\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__9115\ : InMux
    port map (
            O => \N__43152\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__9114\ : InMux
    port map (
            O => \N__43149\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__9113\ : InMux
    port map (
            O => \N__43146\,
            I => \bfn_15_29_0_\
        );

    \I__9112\ : CascadeMux
    port map (
            O => \N__43143\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\
        );

    \I__9111\ : InMux
    port map (
            O => \N__43140\,
            I => \N__43137\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__43137\,
            I => \N__43134\
        );

    \I__9109\ : Span4Mux_h
    port map (
            O => \N__43134\,
            I => \N__43131\
        );

    \I__9108\ : Odrv4
    port map (
            O => \N__43131\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19\
        );

    \I__9107\ : InMux
    port map (
            O => \N__43128\,
            I => \N__43125\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__43125\,
            I => \N__43122\
        );

    \I__9105\ : Span4Mux_v
    port map (
            O => \N__43122\,
            I => \N__43118\
        );

    \I__9104\ : InMux
    port map (
            O => \N__43121\,
            I => \N__43115\
        );

    \I__9103\ : Odrv4
    port map (
            O => \N__43118\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__43115\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9101\ : InMux
    port map (
            O => \N__43110\,
            I => \N__43107\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__43107\,
            I => \N__43104\
        );

    \I__9099\ : Span4Mux_v
    port map (
            O => \N__43104\,
            I => \N__43101\
        );

    \I__9098\ : Span4Mux_v
    port map (
            O => \N__43101\,
            I => \N__43097\
        );

    \I__9097\ : InMux
    port map (
            O => \N__43100\,
            I => \N__43094\
        );

    \I__9096\ : Odrv4
    port map (
            O => \N__43097\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__43094\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9094\ : CascadeMux
    port map (
            O => \N__43089\,
            I => \N__43085\
        );

    \I__9093\ : InMux
    port map (
            O => \N__43088\,
            I => \N__43082\
        );

    \I__9092\ : InMux
    port map (
            O => \N__43085\,
            I => \N__43079\
        );

    \I__9091\ : LocalMux
    port map (
            O => \N__43082\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__43079\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__9089\ : InMux
    port map (
            O => \N__43074\,
            I => \N__43071\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__43071\,
            I => \N__43068\
        );

    \I__9087\ : Span4Mux_h
    port map (
            O => \N__43068\,
            I => \N__43064\
        );

    \I__9086\ : InMux
    port map (
            O => \N__43067\,
            I => \N__43061\
        );

    \I__9085\ : Odrv4
    port map (
            O => \N__43064\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9084\ : LocalMux
    port map (
            O => \N__43061\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9083\ : InMux
    port map (
            O => \N__43056\,
            I => \N__43053\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__43053\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\
        );

    \I__9081\ : CascadeMux
    port map (
            O => \N__43050\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_\
        );

    \I__9080\ : InMux
    port map (
            O => \N__43047\,
            I => \N__43044\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__43044\,
            I => \N__43041\
        );

    \I__9078\ : Odrv12
    port map (
            O => \N__43041\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\
        );

    \I__9077\ : InMux
    port map (
            O => \N__43038\,
            I => \N__43035\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__43035\,
            I => \N__43032\
        );

    \I__9075\ : Span4Mux_h
    port map (
            O => \N__43032\,
            I => \N__43028\
        );

    \I__9074\ : InMux
    port map (
            O => \N__43031\,
            I => \N__43025\
        );

    \I__9073\ : Odrv4
    port map (
            O => \N__43028\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__43025\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__9071\ : InMux
    port map (
            O => \N__43020\,
            I => \N__43017\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__43017\,
            I => \N__43014\
        );

    \I__9069\ : Span4Mux_h
    port map (
            O => \N__43014\,
            I => \N__43010\
        );

    \I__9068\ : InMux
    port map (
            O => \N__43013\,
            I => \N__43007\
        );

    \I__9067\ : Odrv4
    port map (
            O => \N__43010\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__43007\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__9065\ : InMux
    port map (
            O => \N__43002\,
            I => \N__42999\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__42999\,
            I => \N__42995\
        );

    \I__9063\ : CascadeMux
    port map (
            O => \N__42998\,
            I => \N__42992\
        );

    \I__9062\ : Span4Mux_h
    port map (
            O => \N__42995\,
            I => \N__42989\
        );

    \I__9061\ : InMux
    port map (
            O => \N__42992\,
            I => \N__42986\
        );

    \I__9060\ : Odrv4
    port map (
            O => \N__42989\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__9059\ : LocalMux
    port map (
            O => \N__42986\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__9058\ : InMux
    port map (
            O => \N__42981\,
            I => \N__42978\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__42978\,
            I => \N__42975\
        );

    \I__9056\ : Span4Mux_h
    port map (
            O => \N__42975\,
            I => \N__42971\
        );

    \I__9055\ : InMux
    port map (
            O => \N__42974\,
            I => \N__42968\
        );

    \I__9054\ : Odrv4
    port map (
            O => \N__42971\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__9053\ : LocalMux
    port map (
            O => \N__42968\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__9052\ : InMux
    port map (
            O => \N__42963\,
            I => \N__42960\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__42960\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\
        );

    \I__9050\ : InMux
    port map (
            O => \N__42957\,
            I => \N__42954\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__42954\,
            I => \N__42951\
        );

    \I__9048\ : Span12Mux_v
    port map (
            O => \N__42951\,
            I => \N__42947\
        );

    \I__9047\ : InMux
    port map (
            O => \N__42950\,
            I => \N__42944\
        );

    \I__9046\ : Odrv12
    port map (
            O => \N__42947\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__42944\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__9044\ : InMux
    port map (
            O => \N__42939\,
            I => \N__42936\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__42936\,
            I => \N__42932\
        );

    \I__9042\ : CascadeMux
    port map (
            O => \N__42935\,
            I => \N__42929\
        );

    \I__9041\ : Span4Mux_v
    port map (
            O => \N__42932\,
            I => \N__42926\
        );

    \I__9040\ : InMux
    port map (
            O => \N__42929\,
            I => \N__42923\
        );

    \I__9039\ : Odrv4
    port map (
            O => \N__42926\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__42923\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__9037\ : InMux
    port map (
            O => \N__42918\,
            I => \N__42915\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__42915\,
            I => \N__42912\
        );

    \I__9035\ : Span4Mux_v
    port map (
            O => \N__42912\,
            I => \N__42909\
        );

    \I__9034\ : Span4Mux_v
    port map (
            O => \N__42909\,
            I => \N__42905\
        );

    \I__9033\ : InMux
    port map (
            O => \N__42908\,
            I => \N__42902\
        );

    \I__9032\ : Odrv4
    port map (
            O => \N__42905\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__42902\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__9030\ : InMux
    port map (
            O => \N__42897\,
            I => \N__42894\
        );

    \I__9029\ : LocalMux
    port map (
            O => \N__42894\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\
        );

    \I__9028\ : InMux
    port map (
            O => \N__42891\,
            I => \N__42888\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__42888\,
            I => \N__42885\
        );

    \I__9026\ : Span12Mux_h
    port map (
            O => \N__42885\,
            I => \N__42882\
        );

    \I__9025\ : Odrv12
    port map (
            O => \N__42882\,
            I => \pwm_generator_inst.O_12\
        );

    \I__9024\ : InMux
    port map (
            O => \N__42879\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__9023\ : InMux
    port map (
            O => \N__42876\,
            I => \N__42873\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__42873\,
            I => \N__42869\
        );

    \I__9021\ : InMux
    port map (
            O => \N__42872\,
            I => \N__42866\
        );

    \I__9020\ : Span4Mux_v
    port map (
            O => \N__42869\,
            I => \N__42863\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__42866\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__9018\ : Odrv4
    port map (
            O => \N__42863\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__9017\ : InMux
    port map (
            O => \N__42858\,
            I => \N__42855\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__42855\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28\
        );

    \I__9015\ : InMux
    port map (
            O => \N__42852\,
            I => \N__42849\
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__42849\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__9013\ : CascadeMux
    port map (
            O => \N__42846\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29_cascade_\
        );

    \I__9012\ : InMux
    port map (
            O => \N__42843\,
            I => \N__42840\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__42840\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29\
        );

    \I__9010\ : InMux
    port map (
            O => \N__42837\,
            I => \N__42834\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__42834\,
            I => \N__42831\
        );

    \I__9008\ : Span4Mux_v
    port map (
            O => \N__42831\,
            I => \N__42827\
        );

    \I__9007\ : InMux
    port map (
            O => \N__42830\,
            I => \N__42824\
        );

    \I__9006\ : Odrv4
    port map (
            O => \N__42827\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__42824\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__9004\ : InMux
    port map (
            O => \N__42819\,
            I => \N__42816\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__42816\,
            I => \N__42813\
        );

    \I__9002\ : Span4Mux_v
    port map (
            O => \N__42813\,
            I => \N__42810\
        );

    \I__9001\ : Odrv4
    port map (
            O => \N__42810\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\
        );

    \I__9000\ : InMux
    port map (
            O => \N__42807\,
            I => \N__42804\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__42804\,
            I => \N__42801\
        );

    \I__8998\ : Span4Mux_v
    port map (
            O => \N__42801\,
            I => \N__42798\
        );

    \I__8997\ : Span4Mux_v
    port map (
            O => \N__42798\,
            I => \N__42794\
        );

    \I__8996\ : InMux
    port map (
            O => \N__42797\,
            I => \N__42791\
        );

    \I__8995\ : Odrv4
    port map (
            O => \N__42794\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__8994\ : LocalMux
    port map (
            O => \N__42791\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__8993\ : InMux
    port map (
            O => \N__42786\,
            I => \N__42783\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__42783\,
            I => \N__42780\
        );

    \I__8991\ : Span4Mux_h
    port map (
            O => \N__42780\,
            I => \N__42776\
        );

    \I__8990\ : InMux
    port map (
            O => \N__42779\,
            I => \N__42773\
        );

    \I__8989\ : Odrv4
    port map (
            O => \N__42776\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__42773\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__8987\ : InMux
    port map (
            O => \N__42768\,
            I => \N__42765\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__42765\,
            I => \N__42762\
        );

    \I__8985\ : Span4Mux_v
    port map (
            O => \N__42762\,
            I => \N__42758\
        );

    \I__8984\ : CascadeMux
    port map (
            O => \N__42761\,
            I => \N__42755\
        );

    \I__8983\ : Span4Mux_v
    port map (
            O => \N__42758\,
            I => \N__42752\
        );

    \I__8982\ : InMux
    port map (
            O => \N__42755\,
            I => \N__42749\
        );

    \I__8981\ : Odrv4
    port map (
            O => \N__42752\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__42749\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__8979\ : InMux
    port map (
            O => \N__42744\,
            I => \N__42741\
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__42741\,
            I => \N__42738\
        );

    \I__8977\ : Span4Mux_v
    port map (
            O => \N__42738\,
            I => \N__42735\
        );

    \I__8976\ : Span4Mux_v
    port map (
            O => \N__42735\,
            I => \N__42731\
        );

    \I__8975\ : InMux
    port map (
            O => \N__42734\,
            I => \N__42728\
        );

    \I__8974\ : Odrv4
    port map (
            O => \N__42731\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__42728\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__8972\ : InMux
    port map (
            O => \N__42723\,
            I => \N__42720\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__42720\,
            I => \N__42717\
        );

    \I__8970\ : Span4Mux_h
    port map (
            O => \N__42717\,
            I => \N__42713\
        );

    \I__8969\ : InMux
    port map (
            O => \N__42716\,
            I => \N__42710\
        );

    \I__8968\ : Odrv4
    port map (
            O => \N__42713\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__42710\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__8966\ : CascadeMux
    port map (
            O => \N__42705\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\
        );

    \I__8965\ : InMux
    port map (
            O => \N__42702\,
            I => \N__42699\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__42699\,
            I => \N__42696\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__42696\,
            I => \N__42693\
        );

    \I__8962\ : Span4Mux_v
    port map (
            O => \N__42693\,
            I => \N__42689\
        );

    \I__8961\ : InMux
    port map (
            O => \N__42692\,
            I => \N__42686\
        );

    \I__8960\ : Odrv4
    port map (
            O => \N__42689\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__42686\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__8958\ : InMux
    port map (
            O => \N__42681\,
            I => \N__42678\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__42678\,
            I => \N__42675\
        );

    \I__8956\ : Odrv12
    port map (
            O => \N__42675\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\
        );

    \I__8955\ : InMux
    port map (
            O => \N__42672\,
            I => \N__42669\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__42669\,
            I => \N__42666\
        );

    \I__8953\ : Span4Mux_h
    port map (
            O => \N__42666\,
            I => \N__42663\
        );

    \I__8952\ : Sp12to4
    port map (
            O => \N__42663\,
            I => \N__42659\
        );

    \I__8951\ : InMux
    port map (
            O => \N__42662\,
            I => \N__42656\
        );

    \I__8950\ : Odrv12
    port map (
            O => \N__42659\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__42656\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__8948\ : InMux
    port map (
            O => \N__42651\,
            I => \N__42648\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__42648\,
            I => \N__42645\
        );

    \I__8946\ : Span4Mux_h
    port map (
            O => \N__42645\,
            I => \N__42642\
        );

    \I__8945\ : Span4Mux_v
    port map (
            O => \N__42642\,
            I => \N__42638\
        );

    \I__8944\ : InMux
    port map (
            O => \N__42641\,
            I => \N__42635\
        );

    \I__8943\ : Odrv4
    port map (
            O => \N__42638\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__42635\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__8941\ : InMux
    port map (
            O => \N__42630\,
            I => \N__42627\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__42627\,
            I => \N__42624\
        );

    \I__8939\ : Span4Mux_v
    port map (
            O => \N__42624\,
            I => \N__42620\
        );

    \I__8938\ : InMux
    port map (
            O => \N__42623\,
            I => \N__42617\
        );

    \I__8937\ : Odrv4
    port map (
            O => \N__42620\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__42617\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__8935\ : InMux
    port map (
            O => \N__42612\,
            I => \N__42609\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__42609\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__8933\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42603\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__42603\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__8931\ : CascadeMux
    port map (
            O => \N__42600\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\
        );

    \I__8930\ : InMux
    port map (
            O => \N__42597\,
            I => \N__42594\
        );

    \I__8929\ : LocalMux
    port map (
            O => \N__42594\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22\
        );

    \I__8928\ : InMux
    port map (
            O => \N__42591\,
            I => \N__42588\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__42588\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__8926\ : CascadeMux
    port map (
            O => \N__42585\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23_cascade_\
        );

    \I__8925\ : InMux
    port map (
            O => \N__42582\,
            I => \N__42579\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__42579\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23\
        );

    \I__8923\ : InMux
    port map (
            O => \N__42576\,
            I => \N__42570\
        );

    \I__8922\ : InMux
    port map (
            O => \N__42575\,
            I => \N__42570\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__42570\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__8920\ : InMux
    port map (
            O => \N__42567\,
            I => \N__42564\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__42564\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__8918\ : CascadeMux
    port map (
            O => \N__42561\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\
        );

    \I__8917\ : InMux
    port map (
            O => \N__42558\,
            I => \N__42555\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__42555\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30\
        );

    \I__8915\ : InMux
    port map (
            O => \N__42552\,
            I => \N__42549\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__42549\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27\
        );

    \I__8913\ : CascadeMux
    port map (
            O => \N__42546\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\
        );

    \I__8912\ : InMux
    port map (
            O => \N__42543\,
            I => \N__42540\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__42540\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10\
        );

    \I__8910\ : InMux
    port map (
            O => \N__42537\,
            I => \N__42534\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__42534\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__8908\ : CascadeMux
    port map (
            O => \N__42531\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\
        );

    \I__8907\ : InMux
    port map (
            O => \N__42528\,
            I => \N__42525\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__42525\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14\
        );

    \I__8905\ : InMux
    port map (
            O => \N__42522\,
            I => \N__42518\
        );

    \I__8904\ : InMux
    port map (
            O => \N__42521\,
            I => \N__42515\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__42518\,
            I => \N__42512\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__42515\,
            I => \N__42509\
        );

    \I__8901\ : Odrv4
    port map (
            O => \N__42512\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__8900\ : Odrv12
    port map (
            O => \N__42509\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__8899\ : InMux
    port map (
            O => \N__42504\,
            I => \N__42500\
        );

    \I__8898\ : InMux
    port map (
            O => \N__42503\,
            I => \N__42497\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__42500\,
            I => \N__42494\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__42497\,
            I => \N__42491\
        );

    \I__8895\ : Span4Mux_h
    port map (
            O => \N__42494\,
            I => \N__42488\
        );

    \I__8894\ : Odrv4
    port map (
            O => \N__42491\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__8893\ : Odrv4
    port map (
            O => \N__42488\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__8892\ : InMux
    port map (
            O => \N__42483\,
            I => \N__42480\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__42480\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__8890\ : CascadeMux
    port map (
            O => \N__42477\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\
        );

    \I__8889\ : InMux
    port map (
            O => \N__42474\,
            I => \N__42471\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__42471\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18\
        );

    \I__8887\ : InMux
    port map (
            O => \N__42468\,
            I => \N__42465\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__42465\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24\
        );

    \I__8885\ : InMux
    port map (
            O => \N__42462\,
            I => \N__42459\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__42459\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__8883\ : CascadeMux
    port map (
            O => \N__42456\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\
        );

    \I__8882\ : InMux
    port map (
            O => \N__42453\,
            I => \N__42450\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__42450\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25\
        );

    \I__8880\ : CascadeMux
    port map (
            O => \N__42447\,
            I => \N__42444\
        );

    \I__8879\ : InMux
    port map (
            O => \N__42444\,
            I => \N__42441\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__42441\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5\
        );

    \I__8877\ : InMux
    port map (
            O => \N__42438\,
            I => \N__42435\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__42435\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__8875\ : CascadeMux
    port map (
            O => \N__42432\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\
        );

    \I__8874\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42426\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__42426\,
            I => \N__42423\
        );

    \I__8872\ : Span4Mux_v
    port map (
            O => \N__42423\,
            I => \N__42420\
        );

    \I__8871\ : Odrv4
    port map (
            O => \N__42420\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20\
        );

    \I__8870\ : InMux
    port map (
            O => \N__42417\,
            I => \N__42414\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__42414\,
            I => \N__42410\
        );

    \I__8868\ : InMux
    port map (
            O => \N__42413\,
            I => \N__42407\
        );

    \I__8867\ : Span4Mux_h
    port map (
            O => \N__42410\,
            I => \N__42404\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__42407\,
            I => \N__42399\
        );

    \I__8865\ : Span4Mux_h
    port map (
            O => \N__42404\,
            I => \N__42396\
        );

    \I__8864\ : InMux
    port map (
            O => \N__42403\,
            I => \N__42391\
        );

    \I__8863\ : InMux
    port map (
            O => \N__42402\,
            I => \N__42391\
        );

    \I__8862\ : Span4Mux_v
    port map (
            O => \N__42399\,
            I => \N__42388\
        );

    \I__8861\ : Span4Mux_h
    port map (
            O => \N__42396\,
            I => \N__42385\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__42391\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__8859\ : Odrv4
    port map (
            O => \N__42388\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__8858\ : Odrv4
    port map (
            O => \N__42385\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__8857\ : InMux
    port map (
            O => \N__42378\,
            I => \N__42374\
        );

    \I__8856\ : InMux
    port map (
            O => \N__42377\,
            I => \N__42371\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__42374\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__42371\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__8853\ : InMux
    port map (
            O => \N__42366\,
            I => \N__42363\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__42363\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3\
        );

    \I__8851\ : InMux
    port map (
            O => \N__42360\,
            I => \N__42357\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__42357\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__8849\ : CascadeMux
    port map (
            O => \N__42354\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\
        );

    \I__8848\ : InMux
    port map (
            O => \N__42351\,
            I => \N__42348\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__42348\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16\
        );

    \I__8846\ : InMux
    port map (
            O => \N__42345\,
            I => \N__42342\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__42342\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8\
        );

    \I__8844\ : InMux
    port map (
            O => \N__42339\,
            I => \N__42336\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__42336\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__8842\ : InMux
    port map (
            O => \N__42333\,
            I => \N__42330\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__42330\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__8840\ : CascadeMux
    port map (
            O => \N__42327\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7_cascade_\
        );

    \I__8839\ : InMux
    port map (
            O => \N__42324\,
            I => \N__42321\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__42321\,
            I => \N__42318\
        );

    \I__8837\ : Odrv4
    port map (
            O => \N__42318\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7\
        );

    \I__8836\ : InMux
    port map (
            O => \N__42315\,
            I => \N__42309\
        );

    \I__8835\ : InMux
    port map (
            O => \N__42314\,
            I => \N__42309\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__42309\,
            I => \N__42306\
        );

    \I__8833\ : Span4Mux_v
    port map (
            O => \N__42306\,
            I => \N__42303\
        );

    \I__8832\ : Span4Mux_v
    port map (
            O => \N__42303\,
            I => \N__42300\
        );

    \I__8831\ : Odrv4
    port map (
            O => \N__42300\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__8830\ : InMux
    port map (
            O => \N__42297\,
            I => \N__42291\
        );

    \I__8829\ : InMux
    port map (
            O => \N__42296\,
            I => \N__42288\
        );

    \I__8828\ : InMux
    port map (
            O => \N__42295\,
            I => \N__42285\
        );

    \I__8827\ : InMux
    port map (
            O => \N__42294\,
            I => \N__42282\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__42291\,
            I => \N__42277\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__42288\,
            I => \N__42274\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__42285\,
            I => \N__42271\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__42282\,
            I => \N__42268\
        );

    \I__8822\ : InMux
    port map (
            O => \N__42281\,
            I => \N__42265\
        );

    \I__8821\ : InMux
    port map (
            O => \N__42280\,
            I => \N__42262\
        );

    \I__8820\ : Span12Mux_v
    port map (
            O => \N__42277\,
            I => \N__42257\
        );

    \I__8819\ : Span12Mux_v
    port map (
            O => \N__42274\,
            I => \N__42257\
        );

    \I__8818\ : Span4Mux_h
    port map (
            O => \N__42271\,
            I => \N__42254\
        );

    \I__8817\ : Span4Mux_v
    port map (
            O => \N__42268\,
            I => \N__42249\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__42265\,
            I => \N__42249\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__42262\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__8814\ : Odrv12
    port map (
            O => \N__42257\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__8813\ : Odrv4
    port map (
            O => \N__42254\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__8812\ : Odrv4
    port map (
            O => \N__42249\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__8811\ : InMux
    port map (
            O => \N__42240\,
            I => \N__42237\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__42237\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\
        );

    \I__8809\ : InMux
    port map (
            O => \N__42234\,
            I => \N__42231\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__42231\,
            I => \N__42227\
        );

    \I__8807\ : CascadeMux
    port map (
            O => \N__42230\,
            I => \N__42224\
        );

    \I__8806\ : Span4Mux_h
    port map (
            O => \N__42227\,
            I => \N__42220\
        );

    \I__8805\ : InMux
    port map (
            O => \N__42224\,
            I => \N__42217\
        );

    \I__8804\ : InMux
    port map (
            O => \N__42223\,
            I => \N__42214\
        );

    \I__8803\ : Odrv4
    port map (
            O => \N__42220\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__42217\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__42214\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__8800\ : InMux
    port map (
            O => \N__42207\,
            I => \N__42201\
        );

    \I__8799\ : InMux
    port map (
            O => \N__42206\,
            I => \N__42201\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__42201\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__8797\ : InMux
    port map (
            O => \N__42198\,
            I => \N__42194\
        );

    \I__8796\ : InMux
    port map (
            O => \N__42197\,
            I => \N__42191\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__42194\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__42191\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__8793\ : InMux
    port map (
            O => \N__42186\,
            I => \N__42183\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__42183\,
            I => \N__42179\
        );

    \I__8791\ : CascadeMux
    port map (
            O => \N__42182\,
            I => \N__42176\
        );

    \I__8790\ : Span4Mux_h
    port map (
            O => \N__42179\,
            I => \N__42172\
        );

    \I__8789\ : InMux
    port map (
            O => \N__42176\,
            I => \N__42169\
        );

    \I__8788\ : InMux
    port map (
            O => \N__42175\,
            I => \N__42166\
        );

    \I__8787\ : Odrv4
    port map (
            O => \N__42172\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__42169\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__42166\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__8784\ : CEMux
    port map (
            O => \N__42159\,
            I => \N__42154\
        );

    \I__8783\ : CEMux
    port map (
            O => \N__42158\,
            I => \N__42151\
        );

    \I__8782\ : CEMux
    port map (
            O => \N__42157\,
            I => \N__42148\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__42154\,
            I => \N__42144\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__42151\,
            I => \N__42139\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__42148\,
            I => \N__42139\
        );

    \I__8778\ : CEMux
    port map (
            O => \N__42147\,
            I => \N__42136\
        );

    \I__8777\ : Span4Mux_v
    port map (
            O => \N__42144\,
            I => \N__42128\
        );

    \I__8776\ : Span4Mux_v
    port map (
            O => \N__42139\,
            I => \N__42128\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__42136\,
            I => \N__42128\
        );

    \I__8774\ : CEMux
    port map (
            O => \N__42135\,
            I => \N__42125\
        );

    \I__8773\ : Span4Mux_v
    port map (
            O => \N__42128\,
            I => \N__42120\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__42125\,
            I => \N__42120\
        );

    \I__8771\ : Span4Mux_v
    port map (
            O => \N__42120\,
            I => \N__42117\
        );

    \I__8770\ : Odrv4
    port map (
            O => \N__42117\,
            I => \delay_measurement_inst.delay_tr_timer.N_157_i\
        );

    \I__8769\ : InMux
    port map (
            O => \N__42114\,
            I => \N__42108\
        );

    \I__8768\ : InMux
    port map (
            O => \N__42113\,
            I => \N__42108\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__42108\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__8766\ : InMux
    port map (
            O => \N__42105\,
            I => \N__42101\
        );

    \I__8765\ : InMux
    port map (
            O => \N__42104\,
            I => \N__42098\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__42101\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__42098\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__8762\ : InMux
    port map (
            O => \N__42093\,
            I => \N__42087\
        );

    \I__8761\ : InMux
    port map (
            O => \N__42092\,
            I => \N__42087\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__42087\,
            I => \N__42084\
        );

    \I__8759\ : Span4Mux_v
    port map (
            O => \N__42084\,
            I => \N__42081\
        );

    \I__8758\ : Odrv4
    port map (
            O => \N__42081\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__8757\ : InMux
    port map (
            O => \N__42078\,
            I => \N__42075\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__42075\,
            I => \N__42072\
        );

    \I__8755\ : Span4Mux_v
    port map (
            O => \N__42072\,
            I => \N__42069\
        );

    \I__8754\ : Odrv4
    port map (
            O => \N__42069\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13\
        );

    \I__8753\ : InMux
    port map (
            O => \N__42066\,
            I => \N__42063\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__42063\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__8751\ : CascadeMux
    port map (
            O => \N__42060\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21_cascade_\
        );

    \I__8750\ : InMux
    port map (
            O => \N__42057\,
            I => \N__42054\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__42054\,
            I => \N__42051\
        );

    \I__8748\ : Span4Mux_v
    port map (
            O => \N__42051\,
            I => \N__42048\
        );

    \I__8747\ : Odrv4
    port map (
            O => \N__42048\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21\
        );

    \I__8746\ : InMux
    port map (
            O => \N__42045\,
            I => \N__42041\
        );

    \I__8745\ : InMux
    port map (
            O => \N__42044\,
            I => \N__42038\
        );

    \I__8744\ : LocalMux
    port map (
            O => \N__42041\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__42038\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__8742\ : CascadeMux
    port map (
            O => \N__42033\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\
        );

    \I__8741\ : CascadeMux
    port map (
            O => \N__42030\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\
        );

    \I__8740\ : InMux
    port map (
            O => \N__42027\,
            I => \N__42024\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__42024\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__8738\ : CascadeMux
    port map (
            O => \N__42021\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6_cascade_\
        );

    \I__8737\ : CascadeMux
    port map (
            O => \N__42018\,
            I => \N__42015\
        );

    \I__8736\ : InMux
    port map (
            O => \N__42015\,
            I => \N__42012\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__42012\,
            I => \N__42009\
        );

    \I__8734\ : Odrv4
    port map (
            O => \N__42009\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6\
        );

    \I__8733\ : CascadeMux
    port map (
            O => \N__42006\,
            I => \N__42002\
        );

    \I__8732\ : InMux
    port map (
            O => \N__42005\,
            I => \N__41997\
        );

    \I__8731\ : InMux
    port map (
            O => \N__42002\,
            I => \N__41997\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__41997\,
            I => \N__41994\
        );

    \I__8729\ : Span4Mux_v
    port map (
            O => \N__41994\,
            I => \N__41991\
        );

    \I__8728\ : Odrv4
    port map (
            O => \N__41991\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__8727\ : InMux
    port map (
            O => \N__41988\,
            I => \N__41985\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__41985\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__8725\ : CascadeMux
    port map (
            O => \N__41982\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\
        );

    \I__8724\ : InMux
    port map (
            O => \N__41979\,
            I => \N__41976\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__41976\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__8722\ : CascadeMux
    port map (
            O => \N__41973\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12_cascade_\
        );

    \I__8721\ : InMux
    port map (
            O => \N__41970\,
            I => \N__41967\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__41967\,
            I => \N__41964\
        );

    \I__8719\ : Span4Mux_h
    port map (
            O => \N__41964\,
            I => \N__41961\
        );

    \I__8718\ : Span4Mux_v
    port map (
            O => \N__41961\,
            I => \N__41958\
        );

    \I__8717\ : Odrv4
    port map (
            O => \N__41958\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12\
        );

    \I__8716\ : InMux
    port map (
            O => \N__41955\,
            I => \N__41952\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__41952\,
            I => \N__41949\
        );

    \I__8714\ : Span4Mux_v
    port map (
            O => \N__41949\,
            I => \N__41946\
        );

    \I__8713\ : Odrv4
    port map (
            O => \N__41946\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17\
        );

    \I__8712\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41940\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__41940\,
            I => \N__41937\
        );

    \I__8710\ : Span12Mux_h
    port map (
            O => \N__41937\,
            I => \N__41934\
        );

    \I__8709\ : Odrv12
    port map (
            O => \N__41934\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26\
        );

    \I__8708\ : InMux
    port map (
            O => \N__41931\,
            I => \N__41927\
        );

    \I__8707\ : InMux
    port map (
            O => \N__41930\,
            I => \N__41924\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__41927\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__41924\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__8704\ : InMux
    port map (
            O => \N__41919\,
            I => \N__41916\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__41916\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__8702\ : CascadeMux
    port map (
            O => \N__41913\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\
        );

    \I__8701\ : CascadeMux
    port map (
            O => \N__41910\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\
        );

    \I__8700\ : InMux
    port map (
            O => \N__41907\,
            I => \N__41904\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__41904\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__8698\ : CascadeMux
    port map (
            O => \N__41901\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\
        );

    \I__8697\ : InMux
    port map (
            O => \N__41898\,
            I => \N__41895\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__41895\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__8695\ : CascadeMux
    port map (
            O => \N__41892\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\
        );

    \I__8694\ : InMux
    port map (
            O => \N__41889\,
            I => \N__41886\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__41886\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__8692\ : CascadeMux
    port map (
            O => \N__41883\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\
        );

    \I__8691\ : InMux
    port map (
            O => \N__41880\,
            I => \N__41877\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__41877\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__8689\ : CascadeMux
    port map (
            O => \N__41874\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\
        );

    \I__8688\ : InMux
    port map (
            O => \N__41871\,
            I => \N__41868\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__41868\,
            I => \N__41865\
        );

    \I__8686\ : Span4Mux_v
    port map (
            O => \N__41865\,
            I => \N__41862\
        );

    \I__8685\ : Odrv4
    port map (
            O => \N__41862\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11\
        );

    \I__8684\ : CascadeMux
    port map (
            O => \N__41859\,
            I => \N__41856\
        );

    \I__8683\ : InMux
    port map (
            O => \N__41856\,
            I => \N__41853\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__41853\,
            I => \N__41850\
        );

    \I__8681\ : Odrv4
    port map (
            O => \N__41850\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22\
        );

    \I__8680\ : InMux
    port map (
            O => \N__41847\,
            I => \N__41841\
        );

    \I__8679\ : InMux
    port map (
            O => \N__41846\,
            I => \N__41841\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__41841\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_23\
        );

    \I__8677\ : InMux
    port map (
            O => \N__41838\,
            I => \N__41835\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__41835\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt16\
        );

    \I__8675\ : InMux
    port map (
            O => \N__41832\,
            I => \N__41826\
        );

    \I__8674\ : InMux
    port map (
            O => \N__41831\,
            I => \N__41826\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__41826\,
            I => \N__41822\
        );

    \I__8672\ : InMux
    port map (
            O => \N__41825\,
            I => \N__41819\
        );

    \I__8671\ : Span4Mux_v
    port map (
            O => \N__41822\,
            I => \N__41816\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__41819\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_17\
        );

    \I__8669\ : Odrv4
    port map (
            O => \N__41816\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_17\
        );

    \I__8668\ : CascadeMux
    port map (
            O => \N__41811\,
            I => \N__41807\
        );

    \I__8667\ : CascadeMux
    port map (
            O => \N__41810\,
            I => \N__41804\
        );

    \I__8666\ : InMux
    port map (
            O => \N__41807\,
            I => \N__41799\
        );

    \I__8665\ : InMux
    port map (
            O => \N__41804\,
            I => \N__41799\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__41799\,
            I => \N__41795\
        );

    \I__8663\ : InMux
    port map (
            O => \N__41798\,
            I => \N__41792\
        );

    \I__8662\ : Span4Mux_v
    port map (
            O => \N__41795\,
            I => \N__41789\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__41792\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_16\
        );

    \I__8660\ : Odrv4
    port map (
            O => \N__41789\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_16\
        );

    \I__8659\ : CascadeMux
    port map (
            O => \N__41784\,
            I => \N__41781\
        );

    \I__8658\ : InMux
    port map (
            O => \N__41781\,
            I => \N__41778\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__41778\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16\
        );

    \I__8656\ : InMux
    port map (
            O => \N__41775\,
            I => \N__41769\
        );

    \I__8655\ : InMux
    port map (
            O => \N__41774\,
            I => \N__41769\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__41769\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_17\
        );

    \I__8653\ : InMux
    port map (
            O => \N__41766\,
            I => \N__41763\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__41763\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt18\
        );

    \I__8651\ : InMux
    port map (
            O => \N__41760\,
            I => \N__41754\
        );

    \I__8650\ : InMux
    port map (
            O => \N__41759\,
            I => \N__41754\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__41754\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_18\
        );

    \I__8648\ : InMux
    port map (
            O => \N__41751\,
            I => \N__41745\
        );

    \I__8647\ : InMux
    port map (
            O => \N__41750\,
            I => \N__41745\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__41745\,
            I => \N__41741\
        );

    \I__8645\ : InMux
    port map (
            O => \N__41744\,
            I => \N__41738\
        );

    \I__8644\ : Span4Mux_v
    port map (
            O => \N__41741\,
            I => \N__41735\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__41738\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_19\
        );

    \I__8642\ : Odrv4
    port map (
            O => \N__41735\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_19\
        );

    \I__8641\ : CascadeMux
    port map (
            O => \N__41730\,
            I => \N__41726\
        );

    \I__8640\ : CascadeMux
    port map (
            O => \N__41729\,
            I => \N__41723\
        );

    \I__8639\ : InMux
    port map (
            O => \N__41726\,
            I => \N__41718\
        );

    \I__8638\ : InMux
    port map (
            O => \N__41723\,
            I => \N__41718\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__41718\,
            I => \N__41714\
        );

    \I__8636\ : InMux
    port map (
            O => \N__41717\,
            I => \N__41711\
        );

    \I__8635\ : Span4Mux_v
    port map (
            O => \N__41714\,
            I => \N__41708\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__41711\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_18\
        );

    \I__8633\ : Odrv4
    port map (
            O => \N__41708\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_18\
        );

    \I__8632\ : CascadeMux
    port map (
            O => \N__41703\,
            I => \N__41700\
        );

    \I__8631\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41697\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__41697\,
            I => \N__41694\
        );

    \I__8629\ : Odrv4
    port map (
            O => \N__41694\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18\
        );

    \I__8628\ : InMux
    port map (
            O => \N__41691\,
            I => \N__41688\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__41688\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__8626\ : InMux
    port map (
            O => \N__41685\,
            I => \N__41679\
        );

    \I__8625\ : InMux
    port map (
            O => \N__41684\,
            I => \N__41679\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__41679\,
            I => \N__41675\
        );

    \I__8623\ : InMux
    port map (
            O => \N__41678\,
            I => \N__41672\
        );

    \I__8622\ : Span4Mux_h
    port map (
            O => \N__41675\,
            I => \N__41669\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__41672\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_23\
        );

    \I__8620\ : Odrv4
    port map (
            O => \N__41669\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_23\
        );

    \I__8619\ : InMux
    port map (
            O => \N__41664\,
            I => \N__41658\
        );

    \I__8618\ : InMux
    port map (
            O => \N__41663\,
            I => \N__41658\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__41658\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_22\
        );

    \I__8616\ : CascadeMux
    port map (
            O => \N__41655\,
            I => \N__41651\
        );

    \I__8615\ : CascadeMux
    port map (
            O => \N__41654\,
            I => \N__41648\
        );

    \I__8614\ : InMux
    port map (
            O => \N__41651\,
            I => \N__41643\
        );

    \I__8613\ : InMux
    port map (
            O => \N__41648\,
            I => \N__41643\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__41643\,
            I => \N__41639\
        );

    \I__8611\ : InMux
    port map (
            O => \N__41642\,
            I => \N__41636\
        );

    \I__8610\ : Span4Mux_h
    port map (
            O => \N__41639\,
            I => \N__41633\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__41636\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_22\
        );

    \I__8608\ : Odrv4
    port map (
            O => \N__41633\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_22\
        );

    \I__8607\ : CascadeMux
    port map (
            O => \N__41628\,
            I => \N__41625\
        );

    \I__8606\ : InMux
    port map (
            O => \N__41625\,
            I => \N__41622\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__41622\,
            I => \N__41619\
        );

    \I__8604\ : Odrv4
    port map (
            O => \N__41619\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22\
        );

    \I__8603\ : InMux
    port map (
            O => \N__41616\,
            I => \N__41613\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__41613\,
            I => \N__41609\
        );

    \I__8601\ : InMux
    port map (
            O => \N__41612\,
            I => \N__41606\
        );

    \I__8600\ : Span4Mux_h
    port map (
            O => \N__41609\,
            I => \N__41602\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__41606\,
            I => \N__41599\
        );

    \I__8598\ : InMux
    port map (
            O => \N__41605\,
            I => \N__41596\
        );

    \I__8597\ : Span4Mux_v
    port map (
            O => \N__41602\,
            I => \N__41593\
        );

    \I__8596\ : Span12Mux_v
    port map (
            O => \N__41599\,
            I => \N__41590\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__41596\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_25\
        );

    \I__8594\ : Odrv4
    port map (
            O => \N__41593\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_25\
        );

    \I__8593\ : Odrv12
    port map (
            O => \N__41590\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_25\
        );

    \I__8592\ : CascadeMux
    port map (
            O => \N__41583\,
            I => \N__41579\
        );

    \I__8591\ : CascadeMux
    port map (
            O => \N__41582\,
            I => \N__41576\
        );

    \I__8590\ : InMux
    port map (
            O => \N__41579\,
            I => \N__41573\
        );

    \I__8589\ : InMux
    port map (
            O => \N__41576\,
            I => \N__41570\
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__41573\,
            I => \N__41565\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__41570\,
            I => \N__41565\
        );

    \I__8586\ : Span4Mux_h
    port map (
            O => \N__41565\,
            I => \N__41561\
        );

    \I__8585\ : InMux
    port map (
            O => \N__41564\,
            I => \N__41558\
        );

    \I__8584\ : Span4Mux_v
    port map (
            O => \N__41561\,
            I => \N__41555\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__41558\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_24\
        );

    \I__8582\ : Odrv4
    port map (
            O => \N__41555\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_24\
        );

    \I__8581\ : CascadeMux
    port map (
            O => \N__41550\,
            I => \N__41547\
        );

    \I__8580\ : InMux
    port map (
            O => \N__41547\,
            I => \N__41544\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__41544\,
            I => \N__41541\
        );

    \I__8578\ : Span4Mux_v
    port map (
            O => \N__41541\,
            I => \N__41538\
        );

    \I__8577\ : Odrv4
    port map (
            O => \N__41538\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt24\
        );

    \I__8576\ : InMux
    port map (
            O => \N__41535\,
            I => \N__41532\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__41532\,
            I => \N__41529\
        );

    \I__8574\ : Span4Mux_h
    port map (
            O => \N__41529\,
            I => \N__41526\
        );

    \I__8573\ : Odrv4
    port map (
            O => \N__41526\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt20\
        );

    \I__8572\ : InMux
    port map (
            O => \N__41523\,
            I => \N__41517\
        );

    \I__8571\ : InMux
    port map (
            O => \N__41522\,
            I => \N__41517\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__41517\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_20\
        );

    \I__8569\ : CascadeMux
    port map (
            O => \N__41514\,
            I => \N__41510\
        );

    \I__8568\ : CascadeMux
    port map (
            O => \N__41513\,
            I => \N__41507\
        );

    \I__8567\ : InMux
    port map (
            O => \N__41510\,
            I => \N__41502\
        );

    \I__8566\ : InMux
    port map (
            O => \N__41507\,
            I => \N__41502\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__41502\,
            I => \N__41498\
        );

    \I__8564\ : InMux
    port map (
            O => \N__41501\,
            I => \N__41495\
        );

    \I__8563\ : Span4Mux_v
    port map (
            O => \N__41498\,
            I => \N__41492\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__41495\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_21\
        );

    \I__8561\ : Odrv4
    port map (
            O => \N__41492\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_21\
        );

    \I__8560\ : InMux
    port map (
            O => \N__41487\,
            I => \N__41481\
        );

    \I__8559\ : InMux
    port map (
            O => \N__41486\,
            I => \N__41481\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__41481\,
            I => \N__41477\
        );

    \I__8557\ : InMux
    port map (
            O => \N__41480\,
            I => \N__41474\
        );

    \I__8556\ : Span4Mux_v
    port map (
            O => \N__41477\,
            I => \N__41471\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__41474\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_20\
        );

    \I__8554\ : Odrv4
    port map (
            O => \N__41471\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_20\
        );

    \I__8553\ : CascadeMux
    port map (
            O => \N__41466\,
            I => \N__41463\
        );

    \I__8552\ : InMux
    port map (
            O => \N__41463\,
            I => \N__41460\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__41460\,
            I => \N__41457\
        );

    \I__8550\ : Odrv4
    port map (
            O => \N__41457\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20\
        );

    \I__8549\ : InMux
    port map (
            O => \N__41454\,
            I => \N__41451\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__41451\,
            I => \N__41448\
        );

    \I__8547\ : Span4Mux_h
    port map (
            O => \N__41448\,
            I => \N__41445\
        );

    \I__8546\ : Odrv4
    port map (
            O => \N__41445\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt22\
        );

    \I__8545\ : InMux
    port map (
            O => \N__41442\,
            I => \N__41436\
        );

    \I__8544\ : InMux
    port map (
            O => \N__41441\,
            I => \N__41436\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__41436\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_22\
        );

    \I__8542\ : InMux
    port map (
            O => \N__41433\,
            I => \N__41427\
        );

    \I__8541\ : InMux
    port map (
            O => \N__41432\,
            I => \N__41427\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__41427\,
            I => \N__41423\
        );

    \I__8539\ : InMux
    port map (
            O => \N__41426\,
            I => \N__41420\
        );

    \I__8538\ : Span4Mux_v
    port map (
            O => \N__41423\,
            I => \N__41417\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__41420\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_23\
        );

    \I__8536\ : Odrv4
    port map (
            O => \N__41417\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_23\
        );

    \I__8535\ : CascadeMux
    port map (
            O => \N__41412\,
            I => \N__41408\
        );

    \I__8534\ : CascadeMux
    port map (
            O => \N__41411\,
            I => \N__41405\
        );

    \I__8533\ : InMux
    port map (
            O => \N__41408\,
            I => \N__41400\
        );

    \I__8532\ : InMux
    port map (
            O => \N__41405\,
            I => \N__41400\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__41400\,
            I => \N__41396\
        );

    \I__8530\ : InMux
    port map (
            O => \N__41399\,
            I => \N__41393\
        );

    \I__8529\ : Span12Mux_s11_h
    port map (
            O => \N__41396\,
            I => \N__41390\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__41393\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_22\
        );

    \I__8527\ : Odrv12
    port map (
            O => \N__41390\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_22\
        );

    \I__8526\ : InMux
    port map (
            O => \N__41385\,
            I => \N__41382\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__41382\,
            I => \N__41379\
        );

    \I__8524\ : Span4Mux_v
    port map (
            O => \N__41379\,
            I => \N__41376\
        );

    \I__8523\ : Odrv4
    port map (
            O => \N__41376\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_12\
        );

    \I__8522\ : InMux
    port map (
            O => \N__41373\,
            I => \N__41370\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__41370\,
            I => \N__41367\
        );

    \I__8520\ : Odrv4
    port map (
            O => \N__41367\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ1Z_1\
        );

    \I__8519\ : InMux
    port map (
            O => \N__41364\,
            I => \N__41361\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__41361\,
            I => \N__41358\
        );

    \I__8517\ : Span4Mux_v
    port map (
            O => \N__41358\,
            I => \N__41355\
        );

    \I__8516\ : Odrv4
    port map (
            O => \N__41355\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_11\
        );

    \I__8515\ : InMux
    port map (
            O => \N__41352\,
            I => \N__41349\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__41349\,
            I => \N__41346\
        );

    \I__8513\ : Odrv4
    port map (
            O => \N__41346\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_2\
        );

    \I__8512\ : CascadeMux
    port map (
            O => \N__41343\,
            I => \N__41340\
        );

    \I__8511\ : InMux
    port map (
            O => \N__41340\,
            I => \N__41337\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__41337\,
            I => \N__41334\
        );

    \I__8509\ : Odrv12
    port map (
            O => \N__41334\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt20\
        );

    \I__8508\ : InMux
    port map (
            O => \N__41331\,
            I => \N__41325\
        );

    \I__8507\ : InMux
    port map (
            O => \N__41330\,
            I => \N__41325\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__41325\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_20\
        );

    \I__8505\ : InMux
    port map (
            O => \N__41322\,
            I => \N__41316\
        );

    \I__8504\ : InMux
    port map (
            O => \N__41321\,
            I => \N__41316\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__41316\,
            I => \N__41312\
        );

    \I__8502\ : InMux
    port map (
            O => \N__41315\,
            I => \N__41309\
        );

    \I__8501\ : Span4Mux_v
    port map (
            O => \N__41312\,
            I => \N__41306\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__41309\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_21\
        );

    \I__8499\ : Odrv4
    port map (
            O => \N__41306\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_21\
        );

    \I__8498\ : CascadeMux
    port map (
            O => \N__41301\,
            I => \N__41297\
        );

    \I__8497\ : CascadeMux
    port map (
            O => \N__41300\,
            I => \N__41294\
        );

    \I__8496\ : InMux
    port map (
            O => \N__41297\,
            I => \N__41289\
        );

    \I__8495\ : InMux
    port map (
            O => \N__41294\,
            I => \N__41289\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__41289\,
            I => \N__41285\
        );

    \I__8493\ : InMux
    port map (
            O => \N__41288\,
            I => \N__41282\
        );

    \I__8492\ : Span4Mux_v
    port map (
            O => \N__41285\,
            I => \N__41279\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__41282\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_20\
        );

    \I__8490\ : Odrv4
    port map (
            O => \N__41279\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_20\
        );

    \I__8489\ : InMux
    port map (
            O => \N__41274\,
            I => \N__41271\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__41271\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20\
        );

    \I__8487\ : InMux
    port map (
            O => \N__41268\,
            I => \N__41262\
        );

    \I__8486\ : InMux
    port map (
            O => \N__41267\,
            I => \N__41262\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__41262\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_21\
        );

    \I__8484\ : InMux
    port map (
            O => \N__41259\,
            I => \N__41256\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__41256\,
            I => \N__41253\
        );

    \I__8482\ : Odrv4
    port map (
            O => \N__41253\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt22\
        );

    \I__8481\ : IoInMux
    port map (
            O => \N__41250\,
            I => \N__41247\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__41247\,
            I => \N__41244\
        );

    \I__8479\ : Span4Mux_s1_v
    port map (
            O => \N__41244\,
            I => \N__41239\
        );

    \I__8478\ : InMux
    port map (
            O => \N__41243\,
            I => \N__41234\
        );

    \I__8477\ : InMux
    port map (
            O => \N__41242\,
            I => \N__41234\
        );

    \I__8476\ : Odrv4
    port map (
            O => \N__41239\,
            I => s1_phy_c
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__41234\,
            I => s1_phy_c
        );

    \I__8474\ : InMux
    port map (
            O => \N__41229\,
            I => \N__41224\
        );

    \I__8473\ : InMux
    port map (
            O => \N__41228\,
            I => \N__41219\
        );

    \I__8472\ : InMux
    port map (
            O => \N__41227\,
            I => \N__41219\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__41224\,
            I => \N__41212\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__41219\,
            I => \N__41212\
        );

    \I__8469\ : CascadeMux
    port map (
            O => \N__41218\,
            I => \N__41208\
        );

    \I__8468\ : InMux
    port map (
            O => \N__41217\,
            I => \N__41205\
        );

    \I__8467\ : Span4Mux_s3_v
    port map (
            O => \N__41212\,
            I => \N__41202\
        );

    \I__8466\ : CascadeMux
    port map (
            O => \N__41211\,
            I => \N__41199\
        );

    \I__8465\ : InMux
    port map (
            O => \N__41208\,
            I => \N__41196\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__41205\,
            I => \N__41193\
        );

    \I__8463\ : Span4Mux_v
    port map (
            O => \N__41202\,
            I => \N__41190\
        );

    \I__8462\ : InMux
    port map (
            O => \N__41199\,
            I => \N__41187\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__41196\,
            I => \N__41182\
        );

    \I__8460\ : Span4Mux_h
    port map (
            O => \N__41193\,
            I => \N__41182\
        );

    \I__8459\ : Span4Mux_v
    port map (
            O => \N__41190\,
            I => \N__41179\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__41187\,
            I => state_3
        );

    \I__8457\ : Odrv4
    port map (
            O => \N__41182\,
            I => state_3
        );

    \I__8456\ : Odrv4
    port map (
            O => \N__41179\,
            I => state_3
        );

    \I__8455\ : CascadeMux
    port map (
            O => \N__41172\,
            I => \N__41166\
        );

    \I__8454\ : InMux
    port map (
            O => \N__41171\,
            I => \N__41163\
        );

    \I__8453\ : InMux
    port map (
            O => \N__41170\,
            I => \N__41156\
        );

    \I__8452\ : InMux
    port map (
            O => \N__41169\,
            I => \N__41156\
        );

    \I__8451\ : InMux
    port map (
            O => \N__41166\,
            I => \N__41156\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__41163\,
            I => \N__41153\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__41156\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__8448\ : Odrv4
    port map (
            O => \N__41153\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__8447\ : CascadeMux
    port map (
            O => \N__41148\,
            I => \N__41145\
        );

    \I__8446\ : InMux
    port map (
            O => \N__41145\,
            I => \N__41142\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__41142\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_0\
        );

    \I__8444\ : CascadeMux
    port map (
            O => \N__41139\,
            I => \N__41136\
        );

    \I__8443\ : InMux
    port map (
            O => \N__41136\,
            I => \N__41133\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__41133\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_3\
        );

    \I__8441\ : CascadeMux
    port map (
            O => \N__41130\,
            I => \N__41127\
        );

    \I__8440\ : InMux
    port map (
            O => \N__41127\,
            I => \N__41124\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__41124\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_4\
        );

    \I__8438\ : CascadeMux
    port map (
            O => \N__41121\,
            I => \N__41118\
        );

    \I__8437\ : InMux
    port map (
            O => \N__41118\,
            I => \N__41115\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__41115\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_1\
        );

    \I__8435\ : CascadeMux
    port map (
            O => \N__41112\,
            I => \N__41109\
        );

    \I__8434\ : InMux
    port map (
            O => \N__41109\,
            I => \N__41106\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__41106\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_2\
        );

    \I__8432\ : InMux
    port map (
            O => \N__41103\,
            I => \N__41100\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__41100\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_6\
        );

    \I__8430\ : InMux
    port map (
            O => \N__41097\,
            I => \N__41094\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__41094\,
            I => \N__41091\
        );

    \I__8428\ : Span4Mux_v
    port map (
            O => \N__41091\,
            I => \N__41088\
        );

    \I__8427\ : Odrv4
    port map (
            O => \N__41088\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_6\
        );

    \I__8426\ : InMux
    port map (
            O => \N__41085\,
            I => \N__41082\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__41082\,
            I => \N__41079\
        );

    \I__8424\ : Span4Mux_v
    port map (
            O => \N__41079\,
            I => \N__41076\
        );

    \I__8423\ : Odrv4
    port map (
            O => \N__41076\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_8\
        );

    \I__8422\ : CascadeMux
    port map (
            O => \N__41073\,
            I => \N__41070\
        );

    \I__8421\ : InMux
    port map (
            O => \N__41070\,
            I => \N__41065\
        );

    \I__8420\ : InMux
    port map (
            O => \N__41069\,
            I => \N__41062\
        );

    \I__8419\ : InMux
    port map (
            O => \N__41068\,
            I => \N__41059\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__41065\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__41062\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__41059\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__8415\ : InMux
    port map (
            O => \N__41052\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__8414\ : CascadeMux
    port map (
            O => \N__41049\,
            I => \N__41046\
        );

    \I__8413\ : InMux
    port map (
            O => \N__41046\,
            I => \N__41041\
        );

    \I__8412\ : InMux
    port map (
            O => \N__41045\,
            I => \N__41038\
        );

    \I__8411\ : InMux
    port map (
            O => \N__41044\,
            I => \N__41035\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__41041\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__41038\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__41035\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__8407\ : InMux
    port map (
            O => \N__41028\,
            I => \bfn_14_27_0_\
        );

    \I__8406\ : InMux
    port map (
            O => \N__41025\,
            I => \N__41020\
        );

    \I__8405\ : InMux
    port map (
            O => \N__41024\,
            I => \N__41017\
        );

    \I__8404\ : InMux
    port map (
            O => \N__41023\,
            I => \N__41014\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__41020\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__41017\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__41014\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__8400\ : InMux
    port map (
            O => \N__41007\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__8399\ : InMux
    port map (
            O => \N__41004\,
            I => \N__41000\
        );

    \I__8398\ : InMux
    port map (
            O => \N__41003\,
            I => \N__40997\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__41000\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__40997\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__8395\ : CascadeMux
    port map (
            O => \N__40992\,
            I => \N__40989\
        );

    \I__8394\ : InMux
    port map (
            O => \N__40989\,
            I => \N__40984\
        );

    \I__8393\ : InMux
    port map (
            O => \N__40988\,
            I => \N__40981\
        );

    \I__8392\ : InMux
    port map (
            O => \N__40987\,
            I => \N__40978\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__40984\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__40981\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__40978\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__8388\ : InMux
    port map (
            O => \N__40971\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__8387\ : InMux
    port map (
            O => \N__40968\,
            I => \N__40964\
        );

    \I__8386\ : InMux
    port map (
            O => \N__40967\,
            I => \N__40961\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__40964\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__40961\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__8383\ : CascadeMux
    port map (
            O => \N__40956\,
            I => \N__40951\
        );

    \I__8382\ : CascadeMux
    port map (
            O => \N__40955\,
            I => \N__40948\
        );

    \I__8381\ : InMux
    port map (
            O => \N__40954\,
            I => \N__40945\
        );

    \I__8380\ : InMux
    port map (
            O => \N__40951\,
            I => \N__40940\
        );

    \I__8379\ : InMux
    port map (
            O => \N__40948\,
            I => \N__40940\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__40945\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__40940\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__8376\ : InMux
    port map (
            O => \N__40935\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__8375\ : InMux
    port map (
            O => \N__40932\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__8374\ : InMux
    port map (
            O => \N__40929\,
            I => \N__40926\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__40926\,
            I => \N__40922\
        );

    \I__8372\ : InMux
    port map (
            O => \N__40925\,
            I => \N__40918\
        );

    \I__8371\ : Span4Mux_v
    port map (
            O => \N__40922\,
            I => \N__40915\
        );

    \I__8370\ : InMux
    port map (
            O => \N__40921\,
            I => \N__40911\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__40918\,
            I => \N__40908\
        );

    \I__8368\ : Span4Mux_h
    port map (
            O => \N__40915\,
            I => \N__40905\
        );

    \I__8367\ : InMux
    port map (
            O => \N__40914\,
            I => \N__40902\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__40911\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__8365\ : Odrv12
    port map (
            O => \N__40908\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__8364\ : Odrv4
    port map (
            O => \N__40905\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__40902\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__8362\ : InMux
    port map (
            O => \N__40893\,
            I => \N__40888\
        );

    \I__8361\ : InMux
    port map (
            O => \N__40892\,
            I => \N__40882\
        );

    \I__8360\ : InMux
    port map (
            O => \N__40891\,
            I => \N__40882\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__40888\,
            I => \N__40879\
        );

    \I__8358\ : InMux
    port map (
            O => \N__40887\,
            I => \N__40876\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__40882\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__8356\ : Odrv4
    port map (
            O => \N__40879\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__40876\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__8354\ : CascadeMux
    port map (
            O => \N__40869\,
            I => \N__40866\
        );

    \I__8353\ : InMux
    port map (
            O => \N__40866\,
            I => \N__40861\
        );

    \I__8352\ : InMux
    port map (
            O => \N__40865\,
            I => \N__40858\
        );

    \I__8351\ : InMux
    port map (
            O => \N__40864\,
            I => \N__40855\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__40861\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__40858\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__40855\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__8347\ : InMux
    port map (
            O => \N__40848\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__8346\ : CascadeMux
    port map (
            O => \N__40845\,
            I => \N__40842\
        );

    \I__8345\ : InMux
    port map (
            O => \N__40842\,
            I => \N__40837\
        );

    \I__8344\ : InMux
    port map (
            O => \N__40841\,
            I => \N__40834\
        );

    \I__8343\ : InMux
    port map (
            O => \N__40840\,
            I => \N__40831\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__40837\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__40834\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__40831\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__8339\ : InMux
    port map (
            O => \N__40824\,
            I => \bfn_14_26_0_\
        );

    \I__8338\ : CascadeMux
    port map (
            O => \N__40821\,
            I => \N__40818\
        );

    \I__8337\ : InMux
    port map (
            O => \N__40818\,
            I => \N__40813\
        );

    \I__8336\ : InMux
    port map (
            O => \N__40817\,
            I => \N__40810\
        );

    \I__8335\ : InMux
    port map (
            O => \N__40816\,
            I => \N__40807\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__40813\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__40810\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__40807\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__8331\ : InMux
    port map (
            O => \N__40800\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__8330\ : InMux
    port map (
            O => \N__40797\,
            I => \N__40792\
        );

    \I__8329\ : InMux
    port map (
            O => \N__40796\,
            I => \N__40787\
        );

    \I__8328\ : InMux
    port map (
            O => \N__40795\,
            I => \N__40787\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__40792\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__40787\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__8325\ : InMux
    port map (
            O => \N__40782\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__8324\ : CascadeMux
    port map (
            O => \N__40779\,
            I => \N__40776\
        );

    \I__8323\ : InMux
    port map (
            O => \N__40776\,
            I => \N__40771\
        );

    \I__8322\ : InMux
    port map (
            O => \N__40775\,
            I => \N__40768\
        );

    \I__8321\ : InMux
    port map (
            O => \N__40774\,
            I => \N__40765\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__40771\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__40768\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__40765\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__8317\ : InMux
    port map (
            O => \N__40758\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__8316\ : CascadeMux
    port map (
            O => \N__40755\,
            I => \N__40750\
        );

    \I__8315\ : CascadeMux
    port map (
            O => \N__40754\,
            I => \N__40747\
        );

    \I__8314\ : InMux
    port map (
            O => \N__40753\,
            I => \N__40744\
        );

    \I__8313\ : InMux
    port map (
            O => \N__40750\,
            I => \N__40739\
        );

    \I__8312\ : InMux
    port map (
            O => \N__40747\,
            I => \N__40739\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__40744\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__40739\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__8309\ : InMux
    port map (
            O => \N__40734\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__8308\ : CascadeMux
    port map (
            O => \N__40731\,
            I => \N__40728\
        );

    \I__8307\ : InMux
    port map (
            O => \N__40728\,
            I => \N__40723\
        );

    \I__8306\ : InMux
    port map (
            O => \N__40727\,
            I => \N__40720\
        );

    \I__8305\ : InMux
    port map (
            O => \N__40726\,
            I => \N__40717\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__40723\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__40720\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__40717\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__8301\ : InMux
    port map (
            O => \N__40710\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__8300\ : CascadeMux
    port map (
            O => \N__40707\,
            I => \N__40704\
        );

    \I__8299\ : InMux
    port map (
            O => \N__40704\,
            I => \N__40699\
        );

    \I__8298\ : InMux
    port map (
            O => \N__40703\,
            I => \N__40696\
        );

    \I__8297\ : InMux
    port map (
            O => \N__40702\,
            I => \N__40693\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__40699\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__40696\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__40693\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__8293\ : InMux
    port map (
            O => \N__40686\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__8292\ : CascadeMux
    port map (
            O => \N__40683\,
            I => \N__40680\
        );

    \I__8291\ : InMux
    port map (
            O => \N__40680\,
            I => \N__40675\
        );

    \I__8290\ : InMux
    port map (
            O => \N__40679\,
            I => \N__40672\
        );

    \I__8289\ : InMux
    port map (
            O => \N__40678\,
            I => \N__40669\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__40675\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__40672\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__40669\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__8285\ : InMux
    port map (
            O => \N__40662\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__8284\ : CascadeMux
    port map (
            O => \N__40659\,
            I => \N__40656\
        );

    \I__8283\ : InMux
    port map (
            O => \N__40656\,
            I => \N__40651\
        );

    \I__8282\ : InMux
    port map (
            O => \N__40655\,
            I => \N__40648\
        );

    \I__8281\ : InMux
    port map (
            O => \N__40654\,
            I => \N__40645\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__40651\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__40648\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__40645\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__8277\ : InMux
    port map (
            O => \N__40638\,
            I => \bfn_14_25_0_\
        );

    \I__8276\ : InMux
    port map (
            O => \N__40635\,
            I => \N__40630\
        );

    \I__8275\ : InMux
    port map (
            O => \N__40634\,
            I => \N__40627\
        );

    \I__8274\ : InMux
    port map (
            O => \N__40633\,
            I => \N__40624\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__40630\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__40627\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__40624\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__8270\ : InMux
    port map (
            O => \N__40617\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__8269\ : CascadeMux
    port map (
            O => \N__40614\,
            I => \N__40611\
        );

    \I__8268\ : InMux
    port map (
            O => \N__40611\,
            I => \N__40606\
        );

    \I__8267\ : InMux
    port map (
            O => \N__40610\,
            I => \N__40603\
        );

    \I__8266\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40600\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__40606\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__40603\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__40600\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__8262\ : InMux
    port map (
            O => \N__40593\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__8261\ : CascadeMux
    port map (
            O => \N__40590\,
            I => \N__40585\
        );

    \I__8260\ : CascadeMux
    port map (
            O => \N__40589\,
            I => \N__40582\
        );

    \I__8259\ : InMux
    port map (
            O => \N__40588\,
            I => \N__40579\
        );

    \I__8258\ : InMux
    port map (
            O => \N__40585\,
            I => \N__40574\
        );

    \I__8257\ : InMux
    port map (
            O => \N__40582\,
            I => \N__40574\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__40579\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__40574\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__8254\ : InMux
    port map (
            O => \N__40569\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__8253\ : CascadeMux
    port map (
            O => \N__40566\,
            I => \N__40563\
        );

    \I__8252\ : InMux
    port map (
            O => \N__40563\,
            I => \N__40558\
        );

    \I__8251\ : InMux
    port map (
            O => \N__40562\,
            I => \N__40555\
        );

    \I__8250\ : InMux
    port map (
            O => \N__40561\,
            I => \N__40552\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__40558\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__40555\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__40552\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__8246\ : InMux
    port map (
            O => \N__40545\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__8245\ : CascadeMux
    port map (
            O => \N__40542\,
            I => \N__40539\
        );

    \I__8244\ : InMux
    port map (
            O => \N__40539\,
            I => \N__40534\
        );

    \I__8243\ : InMux
    port map (
            O => \N__40538\,
            I => \N__40531\
        );

    \I__8242\ : InMux
    port map (
            O => \N__40537\,
            I => \N__40528\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__40534\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__40531\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__40528\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__8238\ : InMux
    port map (
            O => \N__40521\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__8237\ : CascadeMux
    port map (
            O => \N__40518\,
            I => \N__40515\
        );

    \I__8236\ : InMux
    port map (
            O => \N__40515\,
            I => \N__40510\
        );

    \I__8235\ : InMux
    port map (
            O => \N__40514\,
            I => \N__40507\
        );

    \I__8234\ : InMux
    port map (
            O => \N__40513\,
            I => \N__40504\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__40510\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__40507\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__40504\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__8230\ : InMux
    port map (
            O => \N__40497\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__8229\ : InMux
    port map (
            O => \N__40494\,
            I => \N__40490\
        );

    \I__8228\ : InMux
    port map (
            O => \N__40493\,
            I => \N__40487\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__40490\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__40487\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0\
        );

    \I__8225\ : InMux
    port map (
            O => \N__40482\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29\
        );

    \I__8224\ : InMux
    port map (
            O => \N__40479\,
            I => \N__40476\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__40476\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO\
        );

    \I__8222\ : InMux
    port map (
            O => \N__40473\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30\
        );

    \I__8221\ : InMux
    port map (
            O => \N__40470\,
            I => \N__40467\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__40467\,
            I => \N__40464\
        );

    \I__8219\ : Span12Mux_h
    port map (
            O => \N__40464\,
            I => \N__40460\
        );

    \I__8218\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40457\
        );

    \I__8217\ : Span12Mux_v
    port map (
            O => \N__40460\,
            I => \N__40454\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__40457\,
            I => \N__40451\
        );

    \I__8215\ : Odrv12
    port map (
            O => \N__40454\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_28
        );

    \I__8214\ : Odrv4
    port map (
            O => \N__40451\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_28
        );

    \I__8213\ : InMux
    port map (
            O => \N__40446\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__8212\ : InMux
    port map (
            O => \N__40443\,
            I => \N__40438\
        );

    \I__8211\ : InMux
    port map (
            O => \N__40442\,
            I => \N__40433\
        );

    \I__8210\ : InMux
    port map (
            O => \N__40441\,
            I => \N__40433\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__40438\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__40433\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__8207\ : InMux
    port map (
            O => \N__40428\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__8206\ : CascadeMux
    port map (
            O => \N__40425\,
            I => \N__40422\
        );

    \I__8205\ : InMux
    port map (
            O => \N__40422\,
            I => \N__40417\
        );

    \I__8204\ : InMux
    port map (
            O => \N__40421\,
            I => \N__40414\
        );

    \I__8203\ : InMux
    port map (
            O => \N__40420\,
            I => \N__40411\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__40417\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__40414\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__40411\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__8199\ : InMux
    port map (
            O => \N__40404\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__8198\ : CascadeMux
    port map (
            O => \N__40401\,
            I => \N__40396\
        );

    \I__8197\ : CascadeMux
    port map (
            O => \N__40400\,
            I => \N__40393\
        );

    \I__8196\ : InMux
    port map (
            O => \N__40399\,
            I => \N__40390\
        );

    \I__8195\ : InMux
    port map (
            O => \N__40396\,
            I => \N__40385\
        );

    \I__8194\ : InMux
    port map (
            O => \N__40393\,
            I => \N__40385\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__40390\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__40385\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__8191\ : InMux
    port map (
            O => \N__40380\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__40377\,
            I => \N__40374\
        );

    \I__8189\ : InMux
    port map (
            O => \N__40374\,
            I => \N__40369\
        );

    \I__8188\ : InMux
    port map (
            O => \N__40373\,
            I => \N__40366\
        );

    \I__8187\ : InMux
    port map (
            O => \N__40372\,
            I => \N__40363\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__40369\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__40366\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__40363\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__8183\ : InMux
    port map (
            O => \N__40356\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__8182\ : CascadeMux
    port map (
            O => \N__40353\,
            I => \N__40350\
        );

    \I__8181\ : InMux
    port map (
            O => \N__40350\,
            I => \N__40345\
        );

    \I__8180\ : InMux
    port map (
            O => \N__40349\,
            I => \N__40342\
        );

    \I__8179\ : InMux
    port map (
            O => \N__40348\,
            I => \N__40339\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__40345\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__40342\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__40339\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__8175\ : InMux
    port map (
            O => \N__40332\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__8174\ : InMux
    port map (
            O => \N__40329\,
            I => \N__40325\
        );

    \I__8173\ : InMux
    port map (
            O => \N__40328\,
            I => \N__40322\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__40325\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__40322\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0\
        );

    \I__8170\ : InMux
    port map (
            O => \N__40317\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21\
        );

    \I__8169\ : InMux
    port map (
            O => \N__40314\,
            I => \N__40310\
        );

    \I__8168\ : InMux
    port map (
            O => \N__40313\,
            I => \N__40307\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__40310\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__40307\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0\
        );

    \I__8165\ : InMux
    port map (
            O => \N__40302\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22\
        );

    \I__8164\ : InMux
    port map (
            O => \N__40299\,
            I => \N__40295\
        );

    \I__8163\ : InMux
    port map (
            O => \N__40298\,
            I => \N__40292\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__40295\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__40292\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0\
        );

    \I__8160\ : InMux
    port map (
            O => \N__40287\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23\
        );

    \I__8159\ : InMux
    port map (
            O => \N__40284\,
            I => \N__40280\
        );

    \I__8158\ : InMux
    port map (
            O => \N__40283\,
            I => \N__40277\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__40280\,
            I => \N__40274\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__40277\,
            I => \N__40271\
        );

    \I__8155\ : Odrv4
    port map (
            O => \N__40274\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0\
        );

    \I__8154\ : Odrv4
    port map (
            O => \N__40271\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0\
        );

    \I__8153\ : InMux
    port map (
            O => \N__40266\,
            I => \bfn_14_23_0_\
        );

    \I__8152\ : InMux
    port map (
            O => \N__40263\,
            I => \N__40259\
        );

    \I__8151\ : InMux
    port map (
            O => \N__40262\,
            I => \N__40256\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__40259\,
            I => \N__40251\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__40256\,
            I => \N__40251\
        );

    \I__8148\ : Odrv4
    port map (
            O => \N__40251\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0\
        );

    \I__8147\ : InMux
    port map (
            O => \N__40248\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25\
        );

    \I__8146\ : InMux
    port map (
            O => \N__40245\,
            I => \N__40241\
        );

    \I__8145\ : InMux
    port map (
            O => \N__40244\,
            I => \N__40238\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__40241\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__40238\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0\
        );

    \I__8142\ : InMux
    port map (
            O => \N__40233\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26\
        );

    \I__8141\ : InMux
    port map (
            O => \N__40230\,
            I => \N__40226\
        );

    \I__8140\ : InMux
    port map (
            O => \N__40229\,
            I => \N__40223\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__40226\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__40223\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0\
        );

    \I__8137\ : InMux
    port map (
            O => \N__40218\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27\
        );

    \I__8136\ : InMux
    port map (
            O => \N__40215\,
            I => \N__40211\
        );

    \I__8135\ : InMux
    port map (
            O => \N__40214\,
            I => \N__40208\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__40211\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__40208\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0\
        );

    \I__8132\ : InMux
    port map (
            O => \N__40203\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28\
        );

    \I__8131\ : InMux
    port map (
            O => \N__40200\,
            I => \N__40196\
        );

    \I__8130\ : InMux
    port map (
            O => \N__40199\,
            I => \N__40193\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__40196\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__40193\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9\
        );

    \I__8127\ : InMux
    port map (
            O => \N__40188\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12\
        );

    \I__8126\ : InMux
    port map (
            O => \N__40185\,
            I => \N__40181\
        );

    \I__8125\ : InMux
    port map (
            O => \N__40184\,
            I => \N__40178\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__40181\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__40178\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9\
        );

    \I__8122\ : InMux
    port map (
            O => \N__40173\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13\
        );

    \I__8121\ : InMux
    port map (
            O => \N__40170\,
            I => \N__40166\
        );

    \I__8120\ : InMux
    port map (
            O => \N__40169\,
            I => \N__40163\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__40166\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__40163\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9\
        );

    \I__8117\ : InMux
    port map (
            O => \N__40158\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14\
        );

    \I__8116\ : InMux
    port map (
            O => \N__40155\,
            I => \N__40151\
        );

    \I__8115\ : InMux
    port map (
            O => \N__40154\,
            I => \N__40148\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__40151\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__40148\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9\
        );

    \I__8112\ : InMux
    port map (
            O => \N__40143\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15\
        );

    \I__8111\ : InMux
    port map (
            O => \N__40140\,
            I => \N__40136\
        );

    \I__8110\ : InMux
    port map (
            O => \N__40139\,
            I => \N__40133\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__40136\,
            I => \N__40130\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__40133\,
            I => \N__40127\
        );

    \I__8107\ : Odrv4
    port map (
            O => \N__40130\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0\
        );

    \I__8106\ : Odrv4
    port map (
            O => \N__40127\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0\
        );

    \I__8105\ : InMux
    port map (
            O => \N__40122\,
            I => \bfn_14_22_0_\
        );

    \I__8104\ : InMux
    port map (
            O => \N__40119\,
            I => \N__40115\
        );

    \I__8103\ : InMux
    port map (
            O => \N__40118\,
            I => \N__40112\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__40115\,
            I => \N__40107\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__40112\,
            I => \N__40107\
        );

    \I__8100\ : Odrv4
    port map (
            O => \N__40107\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0\
        );

    \I__8099\ : InMux
    port map (
            O => \N__40104\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17\
        );

    \I__8098\ : InMux
    port map (
            O => \N__40101\,
            I => \N__40097\
        );

    \I__8097\ : InMux
    port map (
            O => \N__40100\,
            I => \N__40094\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__40097\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__40094\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0\
        );

    \I__8094\ : InMux
    port map (
            O => \N__40089\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18\
        );

    \I__8093\ : InMux
    port map (
            O => \N__40086\,
            I => \N__40083\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__40083\,
            I => \N__40079\
        );

    \I__8091\ : InMux
    port map (
            O => \N__40082\,
            I => \N__40076\
        );

    \I__8090\ : Span4Mux_h
    port map (
            O => \N__40079\,
            I => \N__40073\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__40076\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0\
        );

    \I__8088\ : Odrv4
    port map (
            O => \N__40073\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0\
        );

    \I__8087\ : InMux
    port map (
            O => \N__40068\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19\
        );

    \I__8086\ : InMux
    port map (
            O => \N__40065\,
            I => \N__40061\
        );

    \I__8085\ : InMux
    port map (
            O => \N__40064\,
            I => \N__40058\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__40061\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__40058\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0\
        );

    \I__8082\ : InMux
    port map (
            O => \N__40053\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20\
        );

    \I__8081\ : InMux
    port map (
            O => \N__40050\,
            I => \N__40046\
        );

    \I__8080\ : InMux
    port map (
            O => \N__40049\,
            I => \N__40043\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__40046\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__40043\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0\
        );

    \I__8077\ : InMux
    port map (
            O => \N__40038\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4\
        );

    \I__8076\ : InMux
    port map (
            O => \N__40035\,
            I => \N__40031\
        );

    \I__8075\ : InMux
    port map (
            O => \N__40034\,
            I => \N__40028\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__40031\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__40028\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0\
        );

    \I__8072\ : InMux
    port map (
            O => \N__40023\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5\
        );

    \I__8071\ : InMux
    port map (
            O => \N__40020\,
            I => \N__40016\
        );

    \I__8070\ : InMux
    port map (
            O => \N__40019\,
            I => \N__40013\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__40016\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__40013\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0\
        );

    \I__8067\ : InMux
    port map (
            O => \N__40008\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6\
        );

    \I__8066\ : InMux
    port map (
            O => \N__40005\,
            I => \N__40001\
        );

    \I__8065\ : InMux
    port map (
            O => \N__40004\,
            I => \N__39998\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__40001\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__39998\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0\
        );

    \I__8062\ : InMux
    port map (
            O => \N__39993\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7\
        );

    \I__8061\ : InMux
    port map (
            O => \N__39990\,
            I => \N__39987\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__39987\,
            I => \N__39984\
        );

    \I__8059\ : Span4Mux_v
    port map (
            O => \N__39984\,
            I => \N__39981\
        );

    \I__8058\ : Odrv4
    port map (
            O => \N__39981\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9\
        );

    \I__8057\ : InMux
    port map (
            O => \N__39978\,
            I => \N__39974\
        );

    \I__8056\ : InMux
    port map (
            O => \N__39977\,
            I => \N__39971\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__39974\,
            I => \N__39968\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__39971\,
            I => \N__39965\
        );

    \I__8053\ : Odrv4
    port map (
            O => \N__39968\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0\
        );

    \I__8052\ : Odrv4
    port map (
            O => \N__39965\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0\
        );

    \I__8051\ : InMux
    port map (
            O => \N__39960\,
            I => \bfn_14_21_0_\
        );

    \I__8050\ : InMux
    port map (
            O => \N__39957\,
            I => \N__39953\
        );

    \I__8049\ : InMux
    port map (
            O => \N__39956\,
            I => \N__39950\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__39953\,
            I => \N__39945\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__39950\,
            I => \N__39945\
        );

    \I__8046\ : Odrv4
    port map (
            O => \N__39945\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0\
        );

    \I__8045\ : InMux
    port map (
            O => \N__39942\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9\
        );

    \I__8044\ : InMux
    port map (
            O => \N__39939\,
            I => \N__39935\
        );

    \I__8043\ : InMux
    port map (
            O => \N__39938\,
            I => \N__39932\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__39935\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__39932\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9\
        );

    \I__8040\ : InMux
    port map (
            O => \N__39927\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10\
        );

    \I__8039\ : InMux
    port map (
            O => \N__39924\,
            I => \N__39920\
        );

    \I__8038\ : InMux
    port map (
            O => \N__39923\,
            I => \N__39917\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__39920\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__39917\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9\
        );

    \I__8035\ : InMux
    port map (
            O => \N__39912\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11\
        );

    \I__8034\ : InMux
    port map (
            O => \N__39909\,
            I => \N__39903\
        );

    \I__8033\ : InMux
    port map (
            O => \N__39908\,
            I => \N__39903\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__39903\,
            I => \N__39899\
        );

    \I__8031\ : InMux
    port map (
            O => \N__39902\,
            I => \N__39896\
        );

    \I__8030\ : Span4Mux_v
    port map (
            O => \N__39899\,
            I => \N__39893\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__39896\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_28\
        );

    \I__8028\ : Odrv4
    port map (
            O => \N__39893\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_28\
        );

    \I__8027\ : InMux
    port map (
            O => \N__39888\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_27\
        );

    \I__8026\ : CascadeMux
    port map (
            O => \N__39885\,
            I => \N__39882\
        );

    \I__8025\ : InMux
    port map (
            O => \N__39882\,
            I => \N__39876\
        );

    \I__8024\ : InMux
    port map (
            O => \N__39881\,
            I => \N__39876\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__39876\,
            I => \N__39872\
        );

    \I__8022\ : InMux
    port map (
            O => \N__39875\,
            I => \N__39869\
        );

    \I__8021\ : Span4Mux_v
    port map (
            O => \N__39872\,
            I => \N__39866\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__39869\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_29\
        );

    \I__8019\ : Odrv4
    port map (
            O => \N__39866\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_29\
        );

    \I__8018\ : InMux
    port map (
            O => \N__39861\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_28\
        );

    \I__8017\ : InMux
    port map (
            O => \N__39858\,
            I => \N__39854\
        );

    \I__8016\ : InMux
    port map (
            O => \N__39857\,
            I => \N__39851\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__39854\,
            I => \N__39845\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__39851\,
            I => \N__39845\
        );

    \I__8013\ : InMux
    port map (
            O => \N__39850\,
            I => \N__39842\
        );

    \I__8012\ : Span4Mux_v
    port map (
            O => \N__39845\,
            I => \N__39839\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__39842\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_30\
        );

    \I__8010\ : Odrv4
    port map (
            O => \N__39839\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_30\
        );

    \I__8009\ : InMux
    port map (
            O => \N__39834\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_29\
        );

    \I__8008\ : InMux
    port map (
            O => \N__39831\,
            I => \N__39791\
        );

    \I__8007\ : InMux
    port map (
            O => \N__39830\,
            I => \N__39791\
        );

    \I__8006\ : InMux
    port map (
            O => \N__39829\,
            I => \N__39791\
        );

    \I__8005\ : InMux
    port map (
            O => \N__39828\,
            I => \N__39791\
        );

    \I__8004\ : InMux
    port map (
            O => \N__39827\,
            I => \N__39782\
        );

    \I__8003\ : InMux
    port map (
            O => \N__39826\,
            I => \N__39782\
        );

    \I__8002\ : InMux
    port map (
            O => \N__39825\,
            I => \N__39782\
        );

    \I__8001\ : InMux
    port map (
            O => \N__39824\,
            I => \N__39782\
        );

    \I__8000\ : InMux
    port map (
            O => \N__39823\,
            I => \N__39773\
        );

    \I__7999\ : InMux
    port map (
            O => \N__39822\,
            I => \N__39773\
        );

    \I__7998\ : InMux
    port map (
            O => \N__39821\,
            I => \N__39773\
        );

    \I__7997\ : InMux
    port map (
            O => \N__39820\,
            I => \N__39773\
        );

    \I__7996\ : InMux
    port map (
            O => \N__39819\,
            I => \N__39764\
        );

    \I__7995\ : InMux
    port map (
            O => \N__39818\,
            I => \N__39764\
        );

    \I__7994\ : InMux
    port map (
            O => \N__39817\,
            I => \N__39764\
        );

    \I__7993\ : InMux
    port map (
            O => \N__39816\,
            I => \N__39764\
        );

    \I__7992\ : InMux
    port map (
            O => \N__39815\,
            I => \N__39755\
        );

    \I__7991\ : InMux
    port map (
            O => \N__39814\,
            I => \N__39755\
        );

    \I__7990\ : InMux
    port map (
            O => \N__39813\,
            I => \N__39755\
        );

    \I__7989\ : InMux
    port map (
            O => \N__39812\,
            I => \N__39755\
        );

    \I__7988\ : InMux
    port map (
            O => \N__39811\,
            I => \N__39746\
        );

    \I__7987\ : InMux
    port map (
            O => \N__39810\,
            I => \N__39746\
        );

    \I__7986\ : InMux
    port map (
            O => \N__39809\,
            I => \N__39746\
        );

    \I__7985\ : InMux
    port map (
            O => \N__39808\,
            I => \N__39746\
        );

    \I__7984\ : InMux
    port map (
            O => \N__39807\,
            I => \N__39737\
        );

    \I__7983\ : InMux
    port map (
            O => \N__39806\,
            I => \N__39737\
        );

    \I__7982\ : InMux
    port map (
            O => \N__39805\,
            I => \N__39737\
        );

    \I__7981\ : InMux
    port map (
            O => \N__39804\,
            I => \N__39737\
        );

    \I__7980\ : InMux
    port map (
            O => \N__39803\,
            I => \N__39728\
        );

    \I__7979\ : InMux
    port map (
            O => \N__39802\,
            I => \N__39728\
        );

    \I__7978\ : InMux
    port map (
            O => \N__39801\,
            I => \N__39728\
        );

    \I__7977\ : InMux
    port map (
            O => \N__39800\,
            I => \N__39728\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__39791\,
            I => \N__39723\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__39782\,
            I => \N__39723\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__39773\,
            I => \phase_controller_inst1.stoper_hc.start_latched_i_0\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__39764\,
            I => \phase_controller_inst1.stoper_hc.start_latched_i_0\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__39755\,
            I => \phase_controller_inst1.stoper_hc.start_latched_i_0\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__39746\,
            I => \phase_controller_inst1.stoper_hc.start_latched_i_0\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__39737\,
            I => \phase_controller_inst1.stoper_hc.start_latched_i_0\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__39728\,
            I => \phase_controller_inst1.stoper_hc.start_latched_i_0\
        );

    \I__7968\ : Odrv4
    port map (
            O => \N__39723\,
            I => \phase_controller_inst1.stoper_hc.start_latched_i_0\
        );

    \I__7967\ : InMux
    port map (
            O => \N__39708\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_30\
        );

    \I__7966\ : InMux
    port map (
            O => \N__39705\,
            I => \N__39701\
        );

    \I__7965\ : InMux
    port map (
            O => \N__39704\,
            I => \N__39698\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__39701\,
            I => \N__39692\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__39698\,
            I => \N__39692\
        );

    \I__7962\ : InMux
    port map (
            O => \N__39697\,
            I => \N__39689\
        );

    \I__7961\ : Span4Mux_v
    port map (
            O => \N__39692\,
            I => \N__39686\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__39689\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_31\
        );

    \I__7959\ : Odrv4
    port map (
            O => \N__39686\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_31\
        );

    \I__7958\ : CEMux
    port map (
            O => \N__39681\,
            I => \N__39676\
        );

    \I__7957\ : CEMux
    port map (
            O => \N__39680\,
            I => \N__39672\
        );

    \I__7956\ : CEMux
    port map (
            O => \N__39679\,
            I => \N__39669\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__39676\,
            I => \N__39666\
        );

    \I__7954\ : CEMux
    port map (
            O => \N__39675\,
            I => \N__39663\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__39672\,
            I => \N__39660\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__39669\,
            I => \N__39657\
        );

    \I__7951\ : Span4Mux_v
    port map (
            O => \N__39666\,
            I => \N__39654\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__39663\,
            I => \N__39649\
        );

    \I__7949\ : Span4Mux_v
    port map (
            O => \N__39660\,
            I => \N__39649\
        );

    \I__7948\ : Span4Mux_v
    port map (
            O => \N__39657\,
            I => \N__39646\
        );

    \I__7947\ : Span4Mux_h
    port map (
            O => \N__39654\,
            I => \N__39641\
        );

    \I__7946\ : Span4Mux_v
    port map (
            O => \N__39649\,
            I => \N__39641\
        );

    \I__7945\ : Span4Mux_h
    port map (
            O => \N__39646\,
            I => \N__39638\
        );

    \I__7944\ : Span4Mux_h
    port map (
            O => \N__39641\,
            I => \N__39635\
        );

    \I__7943\ : Odrv4
    port map (
            O => \N__39638\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7942\ : Odrv4
    port map (
            O => \N__39635\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7941\ : CascadeMux
    port map (
            O => \N__39630\,
            I => \N__39627\
        );

    \I__7940\ : InMux
    port map (
            O => \N__39627\,
            I => \N__39624\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__39624\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1\
        );

    \I__7938\ : InMux
    port map (
            O => \N__39621\,
            I => \N__39618\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__39618\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2\
        );

    \I__7936\ : InMux
    port map (
            O => \N__39615\,
            I => \N__39611\
        );

    \I__7935\ : InMux
    port map (
            O => \N__39614\,
            I => \N__39608\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__39611\,
            I => \N__39605\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__39608\,
            I => \N__39601\
        );

    \I__7932\ : Span4Mux_v
    port map (
            O => \N__39605\,
            I => \N__39598\
        );

    \I__7931\ : CascadeMux
    port map (
            O => \N__39604\,
            I => \N__39595\
        );

    \I__7930\ : Span4Mux_v
    port map (
            O => \N__39601\,
            I => \N__39590\
        );

    \I__7929\ : Span4Mux_v
    port map (
            O => \N__39598\,
            I => \N__39590\
        );

    \I__7928\ : InMux
    port map (
            O => \N__39595\,
            I => \N__39587\
        );

    \I__7927\ : Odrv4
    port map (
            O => \N__39590\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__39587\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1\
        );

    \I__7925\ : InMux
    port map (
            O => \N__39582\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2\
        );

    \I__7924\ : InMux
    port map (
            O => \N__39579\,
            I => \N__39575\
        );

    \I__7923\ : InMux
    port map (
            O => \N__39578\,
            I => \N__39572\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__39575\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__39572\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0\
        );

    \I__7920\ : InMux
    port map (
            O => \N__39567\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3\
        );

    \I__7919\ : InMux
    port map (
            O => \N__39564\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_18\
        );

    \I__7918\ : InMux
    port map (
            O => \N__39561\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_19\
        );

    \I__7917\ : InMux
    port map (
            O => \N__39558\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_20\
        );

    \I__7916\ : InMux
    port map (
            O => \N__39555\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_21\
        );

    \I__7915\ : InMux
    port map (
            O => \N__39552\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_22\
        );

    \I__7914\ : InMux
    port map (
            O => \N__39549\,
            I => \bfn_14_19_0_\
        );

    \I__7913\ : InMux
    port map (
            O => \N__39546\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_24\
        );

    \I__7912\ : InMux
    port map (
            O => \N__39543\,
            I => \N__39536\
        );

    \I__7911\ : InMux
    port map (
            O => \N__39542\,
            I => \N__39536\
        );

    \I__7910\ : InMux
    port map (
            O => \N__39541\,
            I => \N__39533\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__39536\,
            I => \N__39530\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__39533\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_26\
        );

    \I__7907\ : Odrv12
    port map (
            O => \N__39530\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_26\
        );

    \I__7906\ : InMux
    port map (
            O => \N__39525\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_25\
        );

    \I__7905\ : InMux
    port map (
            O => \N__39522\,
            I => \N__39516\
        );

    \I__7904\ : InMux
    port map (
            O => \N__39521\,
            I => \N__39516\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__39516\,
            I => \N__39512\
        );

    \I__7902\ : InMux
    port map (
            O => \N__39515\,
            I => \N__39509\
        );

    \I__7901\ : Span4Mux_h
    port map (
            O => \N__39512\,
            I => \N__39506\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__39509\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_27\
        );

    \I__7899\ : Odrv4
    port map (
            O => \N__39506\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_27\
        );

    \I__7898\ : InMux
    port map (
            O => \N__39501\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_26\
        );

    \I__7897\ : InMux
    port map (
            O => \N__39498\,
            I => \N__39494\
        );

    \I__7896\ : InMux
    port map (
            O => \N__39497\,
            I => \N__39491\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__39494\,
            I => \N__39488\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__39491\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_10\
        );

    \I__7893\ : Odrv12
    port map (
            O => \N__39488\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_10\
        );

    \I__7892\ : InMux
    port map (
            O => \N__39483\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_9\
        );

    \I__7891\ : InMux
    port map (
            O => \N__39480\,
            I => \N__39476\
        );

    \I__7890\ : InMux
    port map (
            O => \N__39479\,
            I => \N__39473\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__39476\,
            I => \N__39470\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__39473\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_11\
        );

    \I__7887\ : Odrv12
    port map (
            O => \N__39470\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_11\
        );

    \I__7886\ : InMux
    port map (
            O => \N__39465\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_10\
        );

    \I__7885\ : InMux
    port map (
            O => \N__39462\,
            I => \N__39459\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__39459\,
            I => \N__39455\
        );

    \I__7883\ : InMux
    port map (
            O => \N__39458\,
            I => \N__39452\
        );

    \I__7882\ : Span4Mux_v
    port map (
            O => \N__39455\,
            I => \N__39449\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__39452\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_12\
        );

    \I__7880\ : Odrv4
    port map (
            O => \N__39449\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_12\
        );

    \I__7879\ : InMux
    port map (
            O => \N__39444\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_11\
        );

    \I__7878\ : InMux
    port map (
            O => \N__39441\,
            I => \N__39437\
        );

    \I__7877\ : InMux
    port map (
            O => \N__39440\,
            I => \N__39434\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__39437\,
            I => \N__39431\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__39434\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_13\
        );

    \I__7874\ : Odrv12
    port map (
            O => \N__39431\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_13\
        );

    \I__7873\ : InMux
    port map (
            O => \N__39426\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_12\
        );

    \I__7872\ : InMux
    port map (
            O => \N__39423\,
            I => \N__39419\
        );

    \I__7871\ : InMux
    port map (
            O => \N__39422\,
            I => \N__39416\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__39419\,
            I => \N__39413\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__39416\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_14\
        );

    \I__7868\ : Odrv12
    port map (
            O => \N__39413\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_14\
        );

    \I__7867\ : InMux
    port map (
            O => \N__39408\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_13\
        );

    \I__7866\ : InMux
    port map (
            O => \N__39405\,
            I => \N__39401\
        );

    \I__7865\ : InMux
    port map (
            O => \N__39404\,
            I => \N__39398\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__39401\,
            I => \N__39395\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__39398\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_15\
        );

    \I__7862\ : Odrv12
    port map (
            O => \N__39395\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_15\
        );

    \I__7861\ : InMux
    port map (
            O => \N__39390\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_14\
        );

    \I__7860\ : InMux
    port map (
            O => \N__39387\,
            I => \bfn_14_18_0_\
        );

    \I__7859\ : InMux
    port map (
            O => \N__39384\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_16\
        );

    \I__7858\ : InMux
    port map (
            O => \N__39381\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_17\
        );

    \I__7857\ : InMux
    port map (
            O => \N__39378\,
            I => \N__39374\
        );

    \I__7856\ : InMux
    port map (
            O => \N__39377\,
            I => \N__39371\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__39374\,
            I => \N__39368\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__39371\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_2\
        );

    \I__7853\ : Odrv12
    port map (
            O => \N__39368\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_2\
        );

    \I__7852\ : InMux
    port map (
            O => \N__39363\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_1\
        );

    \I__7851\ : InMux
    port map (
            O => \N__39360\,
            I => \N__39356\
        );

    \I__7850\ : InMux
    port map (
            O => \N__39359\,
            I => \N__39353\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__39356\,
            I => \N__39350\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__39353\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_3\
        );

    \I__7847\ : Odrv12
    port map (
            O => \N__39350\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_3\
        );

    \I__7846\ : InMux
    port map (
            O => \N__39345\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_2\
        );

    \I__7845\ : InMux
    port map (
            O => \N__39342\,
            I => \N__39338\
        );

    \I__7844\ : InMux
    port map (
            O => \N__39341\,
            I => \N__39335\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__39338\,
            I => \N__39332\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__39335\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_4\
        );

    \I__7841\ : Odrv12
    port map (
            O => \N__39332\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_4\
        );

    \I__7840\ : InMux
    port map (
            O => \N__39327\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_3\
        );

    \I__7839\ : InMux
    port map (
            O => \N__39324\,
            I => \N__39320\
        );

    \I__7838\ : InMux
    port map (
            O => \N__39323\,
            I => \N__39317\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__39320\,
            I => \N__39314\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__39317\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_5\
        );

    \I__7835\ : Odrv12
    port map (
            O => \N__39314\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_5\
        );

    \I__7834\ : InMux
    port map (
            O => \N__39309\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_4\
        );

    \I__7833\ : InMux
    port map (
            O => \N__39306\,
            I => \N__39302\
        );

    \I__7832\ : InMux
    port map (
            O => \N__39305\,
            I => \N__39299\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__39302\,
            I => \N__39296\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__39299\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_6\
        );

    \I__7829\ : Odrv12
    port map (
            O => \N__39296\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_6\
        );

    \I__7828\ : InMux
    port map (
            O => \N__39291\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_5\
        );

    \I__7827\ : InMux
    port map (
            O => \N__39288\,
            I => \N__39284\
        );

    \I__7826\ : InMux
    port map (
            O => \N__39287\,
            I => \N__39281\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__39284\,
            I => \N__39278\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__39281\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_7\
        );

    \I__7823\ : Odrv12
    port map (
            O => \N__39278\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_7\
        );

    \I__7822\ : InMux
    port map (
            O => \N__39273\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_6\
        );

    \I__7821\ : InMux
    port map (
            O => \N__39270\,
            I => \N__39266\
        );

    \I__7820\ : InMux
    port map (
            O => \N__39269\,
            I => \N__39263\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__39266\,
            I => \N__39260\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__39263\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_8\
        );

    \I__7817\ : Odrv12
    port map (
            O => \N__39260\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_8\
        );

    \I__7816\ : InMux
    port map (
            O => \N__39255\,
            I => \bfn_14_17_0_\
        );

    \I__7815\ : InMux
    port map (
            O => \N__39252\,
            I => \N__39248\
        );

    \I__7814\ : InMux
    port map (
            O => \N__39251\,
            I => \N__39245\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__39248\,
            I => \N__39242\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__39245\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_9\
        );

    \I__7811\ : Odrv12
    port map (
            O => \N__39242\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_9\
        );

    \I__7810\ : InMux
    port map (
            O => \N__39237\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_8\
        );

    \I__7809\ : InMux
    port map (
            O => \N__39234\,
            I => \bfn_14_15_0_\
        );

    \I__7808\ : CascadeMux
    port map (
            O => \N__39231\,
            I => \N__39227\
        );

    \I__7807\ : InMux
    port map (
            O => \N__39230\,
            I => \N__39222\
        );

    \I__7806\ : InMux
    port map (
            O => \N__39227\,
            I => \N__39222\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__39222\,
            I => \N__39219\
        );

    \I__7804\ : Span4Mux_h
    port map (
            O => \N__39219\,
            I => \N__39216\
        );

    \I__7803\ : Odrv4
    port map (
            O => \N__39216\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO\
        );

    \I__7802\ : CascadeMux
    port map (
            O => \N__39213\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO_cascade_\
        );

    \I__7801\ : InMux
    port map (
            O => \N__39210\,
            I => \N__39204\
        );

    \I__7800\ : InMux
    port map (
            O => \N__39209\,
            I => \N__39201\
        );

    \I__7799\ : InMux
    port map (
            O => \N__39208\,
            I => \N__39198\
        );

    \I__7798\ : CascadeMux
    port map (
            O => \N__39207\,
            I => \N__39194\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__39204\,
            I => \N__39190\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__39201\,
            I => \N__39187\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__39198\,
            I => \N__39184\
        );

    \I__7794\ : InMux
    port map (
            O => \N__39197\,
            I => \N__39181\
        );

    \I__7793\ : InMux
    port map (
            O => \N__39194\,
            I => \N__39176\
        );

    \I__7792\ : InMux
    port map (
            O => \N__39193\,
            I => \N__39176\
        );

    \I__7791\ : Span4Mux_v
    port map (
            O => \N__39190\,
            I => \N__39173\
        );

    \I__7790\ : Span4Mux_v
    port map (
            O => \N__39187\,
            I => \N__39168\
        );

    \I__7789\ : Span4Mux_v
    port map (
            O => \N__39184\,
            I => \N__39168\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__39181\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__39176\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7786\ : Odrv4
    port map (
            O => \N__39173\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7785\ : Odrv4
    port map (
            O => \N__39168\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7784\ : InMux
    port map (
            O => \N__39159\,
            I => \N__39153\
        );

    \I__7783\ : InMux
    port map (
            O => \N__39158\,
            I => \N__39150\
        );

    \I__7782\ : InMux
    port map (
            O => \N__39157\,
            I => \N__39145\
        );

    \I__7781\ : InMux
    port map (
            O => \N__39156\,
            I => \N__39145\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__39153\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__39150\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__39145\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28\
        );

    \I__7777\ : CascadeMux
    port map (
            O => \N__39138\,
            I => \N__39135\
        );

    \I__7776\ : InMux
    port map (
            O => \N__39135\,
            I => \N__39132\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__39132\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt30\
        );

    \I__7774\ : CascadeMux
    port map (
            O => \N__39129\,
            I => \N__39126\
        );

    \I__7773\ : InMux
    port map (
            O => \N__39126\,
            I => \N__39123\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__39123\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt26\
        );

    \I__7771\ : InMux
    port map (
            O => \N__39120\,
            I => \N__39117\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__39117\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26\
        );

    \I__7769\ : InMux
    port map (
            O => \N__39114\,
            I => \N__39111\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__39111\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__7767\ : CascadeMux
    port map (
            O => \N__39108\,
            I => \elapsed_time_ns_1_RNILK91B_0_9_cascade_\
        );

    \I__7766\ : InMux
    port map (
            O => \N__39105\,
            I => \N__39101\
        );

    \I__7765\ : CascadeMux
    port map (
            O => \N__39104\,
            I => \N__39098\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__39101\,
            I => \N__39095\
        );

    \I__7763\ : InMux
    port map (
            O => \N__39098\,
            I => \N__39092\
        );

    \I__7762\ : Odrv4
    port map (
            O => \N__39095\,
            I => \phase_controller_inst1.stoper_hc.counter\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__39092\,
            I => \phase_controller_inst1.stoper_hc.counter\
        );

    \I__7760\ : InMux
    port map (
            O => \N__39087\,
            I => \N__39083\
        );

    \I__7759\ : InMux
    port map (
            O => \N__39086\,
            I => \N__39080\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__39083\,
            I => \N__39077\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__39080\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_0\
        );

    \I__7756\ : Odrv12
    port map (
            O => \N__39077\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_0\
        );

    \I__7755\ : InMux
    port map (
            O => \N__39072\,
            I => \N__39068\
        );

    \I__7754\ : InMux
    port map (
            O => \N__39071\,
            I => \N__39065\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__39068\,
            I => \N__39062\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__39065\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_1\
        );

    \I__7751\ : Odrv12
    port map (
            O => \N__39062\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_1\
        );

    \I__7750\ : InMux
    port map (
            O => \N__39057\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_0\
        );

    \I__7749\ : CascadeMux
    port map (
            O => \N__39054\,
            I => \N__39051\
        );

    \I__7748\ : InMux
    port map (
            O => \N__39051\,
            I => \N__39048\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__39048\,
            I => \phase_controller_inst1.stoper_hc.counter_i_15\
        );

    \I__7746\ : InMux
    port map (
            O => \N__39045\,
            I => \N__39042\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__39042\,
            I => \N__39039\
        );

    \I__7744\ : Odrv4
    port map (
            O => \N__39039\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24\
        );

    \I__7743\ : InMux
    port map (
            O => \N__39036\,
            I => \N__39033\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__39033\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28\
        );

    \I__7741\ : CascadeMux
    port map (
            O => \N__39030\,
            I => \N__39027\
        );

    \I__7740\ : InMux
    port map (
            O => \N__39027\,
            I => \N__39024\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__39024\,
            I => \N__39021\
        );

    \I__7738\ : Odrv4
    port map (
            O => \N__39021\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt28\
        );

    \I__7737\ : InMux
    port map (
            O => \N__39018\,
            I => \N__39015\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__39015\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30\
        );

    \I__7735\ : CascadeMux
    port map (
            O => \N__39012\,
            I => \N__39009\
        );

    \I__7734\ : InMux
    port map (
            O => \N__39009\,
            I => \N__39006\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__39006\,
            I => \phase_controller_inst1.stoper_hc.counter_i_7\
        );

    \I__7732\ : CascadeMux
    port map (
            O => \N__39003\,
            I => \N__39000\
        );

    \I__7731\ : InMux
    port map (
            O => \N__39000\,
            I => \N__38997\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__38997\,
            I => \phase_controller_inst1.stoper_hc.counter_i_8\
        );

    \I__7729\ : CascadeMux
    port map (
            O => \N__38994\,
            I => \N__38991\
        );

    \I__7728\ : InMux
    port map (
            O => \N__38991\,
            I => \N__38988\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__38988\,
            I => \phase_controller_inst1.stoper_hc.counter_i_9\
        );

    \I__7726\ : CascadeMux
    port map (
            O => \N__38985\,
            I => \N__38982\
        );

    \I__7725\ : InMux
    port map (
            O => \N__38982\,
            I => \N__38979\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__38979\,
            I => \phase_controller_inst1.stoper_hc.counter_i_10\
        );

    \I__7723\ : CascadeMux
    port map (
            O => \N__38976\,
            I => \N__38973\
        );

    \I__7722\ : InMux
    port map (
            O => \N__38973\,
            I => \N__38970\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__38970\,
            I => \N__38967\
        );

    \I__7720\ : Odrv4
    port map (
            O => \N__38967\,
            I => \phase_controller_inst1.stoper_hc.counter_i_11\
        );

    \I__7719\ : CascadeMux
    port map (
            O => \N__38964\,
            I => \N__38961\
        );

    \I__7718\ : InMux
    port map (
            O => \N__38961\,
            I => \N__38958\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__38958\,
            I => \N__38955\
        );

    \I__7716\ : Odrv4
    port map (
            O => \N__38955\,
            I => \phase_controller_inst1.stoper_hc.counter_i_12\
        );

    \I__7715\ : CascadeMux
    port map (
            O => \N__38952\,
            I => \N__38949\
        );

    \I__7714\ : InMux
    port map (
            O => \N__38949\,
            I => \N__38946\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__38946\,
            I => \phase_controller_inst1.stoper_hc.counter_i_13\
        );

    \I__7712\ : CascadeMux
    port map (
            O => \N__38943\,
            I => \N__38940\
        );

    \I__7711\ : InMux
    port map (
            O => \N__38940\,
            I => \N__38937\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__38937\,
            I => \phase_controller_inst1.stoper_hc.counter_i_14\
        );

    \I__7709\ : InMux
    port map (
            O => \N__38934\,
            I => \N__38929\
        );

    \I__7708\ : InMux
    port map (
            O => \N__38933\,
            I => \N__38924\
        );

    \I__7707\ : InMux
    port map (
            O => \N__38932\,
            I => \N__38924\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__38929\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_28\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__38924\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_28\
        );

    \I__7704\ : CascadeMux
    port map (
            O => \N__38919\,
            I => \N__38915\
        );

    \I__7703\ : InMux
    port map (
            O => \N__38918\,
            I => \N__38908\
        );

    \I__7702\ : InMux
    port map (
            O => \N__38915\,
            I => \N__38908\
        );

    \I__7701\ : InMux
    port map (
            O => \N__38914\,
            I => \N__38903\
        );

    \I__7700\ : InMux
    port map (
            O => \N__38913\,
            I => \N__38903\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__38908\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__38903\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28\
        );

    \I__7697\ : InMux
    port map (
            O => \N__38898\,
            I => \N__38893\
        );

    \I__7696\ : InMux
    port map (
            O => \N__38897\,
            I => \N__38888\
        );

    \I__7695\ : InMux
    port map (
            O => \N__38896\,
            I => \N__38888\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__38893\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_29\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__38888\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_29\
        );

    \I__7692\ : InMux
    port map (
            O => \N__38883\,
            I => \N__38880\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__38880\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt28\
        );

    \I__7690\ : InMux
    port map (
            O => \N__38877\,
            I => \N__38874\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__38874\,
            I => \N__38871\
        );

    \I__7688\ : Span4Mux_v
    port map (
            O => \N__38871\,
            I => \N__38868\
        );

    \I__7687\ : Span4Mux_h
    port map (
            O => \N__38868\,
            I => \N__38865\
        );

    \I__7686\ : Odrv4
    port map (
            O => \N__38865\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_0\
        );

    \I__7685\ : CascadeMux
    port map (
            O => \N__38862\,
            I => \N__38859\
        );

    \I__7684\ : InMux
    port map (
            O => \N__38859\,
            I => \N__38856\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__38856\,
            I => \phase_controller_inst1.stoper_hc.counter_i_0\
        );

    \I__7682\ : CascadeMux
    port map (
            O => \N__38853\,
            I => \N__38850\
        );

    \I__7681\ : InMux
    port map (
            O => \N__38850\,
            I => \N__38847\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__38847\,
            I => \phase_controller_inst1.stoper_hc.counter_i_1\
        );

    \I__7679\ : CascadeMux
    port map (
            O => \N__38844\,
            I => \N__38841\
        );

    \I__7678\ : InMux
    port map (
            O => \N__38841\,
            I => \N__38838\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__38838\,
            I => \phase_controller_inst1.stoper_hc.counter_i_2\
        );

    \I__7676\ : CascadeMux
    port map (
            O => \N__38835\,
            I => \N__38832\
        );

    \I__7675\ : InMux
    port map (
            O => \N__38832\,
            I => \N__38829\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__38829\,
            I => \phase_controller_inst1.stoper_hc.counter_i_3\
        );

    \I__7673\ : CascadeMux
    port map (
            O => \N__38826\,
            I => \N__38823\
        );

    \I__7672\ : InMux
    port map (
            O => \N__38823\,
            I => \N__38820\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__38820\,
            I => \N__38817\
        );

    \I__7670\ : Odrv4
    port map (
            O => \N__38817\,
            I => \phase_controller_inst1.stoper_hc.counter_i_4\
        );

    \I__7669\ : CascadeMux
    port map (
            O => \N__38814\,
            I => \N__38811\
        );

    \I__7668\ : InMux
    port map (
            O => \N__38811\,
            I => \N__38808\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__38808\,
            I => \phase_controller_inst1.stoper_hc.counter_i_5\
        );

    \I__7666\ : CascadeMux
    port map (
            O => \N__38805\,
            I => \N__38802\
        );

    \I__7665\ : InMux
    port map (
            O => \N__38802\,
            I => \N__38799\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__38799\,
            I => \phase_controller_inst1.stoper_hc.counter_i_6\
        );

    \I__7663\ : InMux
    port map (
            O => \N__38796\,
            I => \N__38793\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__38793\,
            I => \N__38790\
        );

    \I__7661\ : Odrv4
    port map (
            O => \N__38790\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30\
        );

    \I__7660\ : CascadeMux
    port map (
            O => \N__38787\,
            I => \N__38784\
        );

    \I__7659\ : InMux
    port map (
            O => \N__38784\,
            I => \N__38781\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__38781\,
            I => \N__38778\
        );

    \I__7657\ : Odrv4
    port map (
            O => \N__38778\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt30\
        );

    \I__7656\ : InMux
    port map (
            O => \N__38775\,
            I => \bfn_14_11_0_\
        );

    \I__7655\ : InMux
    port map (
            O => \N__38772\,
            I => \N__38766\
        );

    \I__7654\ : InMux
    port map (
            O => \N__38771\,
            I => \N__38766\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__38766\,
            I => \N__38763\
        );

    \I__7652\ : Span4Mux_v
    port map (
            O => \N__38763\,
            I => \N__38759\
        );

    \I__7651\ : InMux
    port map (
            O => \N__38762\,
            I => \N__38756\
        );

    \I__7650\ : Span4Mux_h
    port map (
            O => \N__38759\,
            I => \N__38753\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__38756\,
            I => \N__38750\
        );

    \I__7648\ : Odrv4
    port map (
            O => \N__38753\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\
        );

    \I__7647\ : Odrv12
    port map (
            O => \N__38750\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\
        );

    \I__7646\ : CascadeMux
    port map (
            O => \N__38745\,
            I => \N__38742\
        );

    \I__7645\ : InMux
    port map (
            O => \N__38742\,
            I => \N__38739\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__38739\,
            I => \N__38736\
        );

    \I__7643\ : Odrv4
    port map (
            O => \N__38736\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28\
        );

    \I__7642\ : InMux
    port map (
            O => \N__38733\,
            I => \N__38729\
        );

    \I__7641\ : InMux
    port map (
            O => \N__38732\,
            I => \N__38726\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__38729\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_10\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__38726\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_10\
        );

    \I__7638\ : CascadeMux
    port map (
            O => \N__38721\,
            I => \N__38718\
        );

    \I__7637\ : InMux
    port map (
            O => \N__38718\,
            I => \N__38715\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__38715\,
            I => \phase_controller_inst2.stoper_hc.counter_i_10\
        );

    \I__7635\ : InMux
    port map (
            O => \N__38712\,
            I => \N__38708\
        );

    \I__7634\ : InMux
    port map (
            O => \N__38711\,
            I => \N__38705\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__38708\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_11\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__38705\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_11\
        );

    \I__7631\ : CascadeMux
    port map (
            O => \N__38700\,
            I => \N__38697\
        );

    \I__7630\ : InMux
    port map (
            O => \N__38697\,
            I => \N__38694\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__38694\,
            I => \phase_controller_inst2.stoper_hc.counter_i_11\
        );

    \I__7628\ : InMux
    port map (
            O => \N__38691\,
            I => \N__38687\
        );

    \I__7627\ : InMux
    port map (
            O => \N__38690\,
            I => \N__38684\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__38687\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_12\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__38684\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_12\
        );

    \I__7624\ : CascadeMux
    port map (
            O => \N__38679\,
            I => \N__38676\
        );

    \I__7623\ : InMux
    port map (
            O => \N__38676\,
            I => \N__38673\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__38673\,
            I => \N__38670\
        );

    \I__7621\ : Odrv4
    port map (
            O => \N__38670\,
            I => \phase_controller_inst2.stoper_hc.counter_i_12\
        );

    \I__7620\ : InMux
    port map (
            O => \N__38667\,
            I => \N__38663\
        );

    \I__7619\ : InMux
    port map (
            O => \N__38666\,
            I => \N__38660\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__38663\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_13\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__38660\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_13\
        );

    \I__7616\ : CascadeMux
    port map (
            O => \N__38655\,
            I => \N__38652\
        );

    \I__7615\ : InMux
    port map (
            O => \N__38652\,
            I => \N__38649\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__38649\,
            I => \phase_controller_inst2.stoper_hc.counter_i_13\
        );

    \I__7613\ : InMux
    port map (
            O => \N__38646\,
            I => \N__38642\
        );

    \I__7612\ : InMux
    port map (
            O => \N__38645\,
            I => \N__38639\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__38642\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_14\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__38639\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_14\
        );

    \I__7609\ : CascadeMux
    port map (
            O => \N__38634\,
            I => \N__38631\
        );

    \I__7608\ : InMux
    port map (
            O => \N__38631\,
            I => \N__38628\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__38628\,
            I => \phase_controller_inst2.stoper_hc.counter_i_14\
        );

    \I__7606\ : InMux
    port map (
            O => \N__38625\,
            I => \N__38621\
        );

    \I__7605\ : InMux
    port map (
            O => \N__38624\,
            I => \N__38618\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__38621\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_15\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__38618\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_15\
        );

    \I__7602\ : CascadeMux
    port map (
            O => \N__38613\,
            I => \N__38610\
        );

    \I__7601\ : InMux
    port map (
            O => \N__38610\,
            I => \N__38607\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__38607\,
            I => \phase_controller_inst2.stoper_hc.counter_i_15\
        );

    \I__7599\ : InMux
    port map (
            O => \N__38604\,
            I => \N__38600\
        );

    \I__7598\ : InMux
    port map (
            O => \N__38603\,
            I => \N__38597\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__38600\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_2\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__38597\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_2\
        );

    \I__7595\ : InMux
    port map (
            O => \N__38592\,
            I => \N__38589\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__38589\,
            I => \phase_controller_inst2.stoper_hc.counter_i_2\
        );

    \I__7593\ : InMux
    port map (
            O => \N__38586\,
            I => \N__38582\
        );

    \I__7592\ : InMux
    port map (
            O => \N__38585\,
            I => \N__38579\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__38582\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_3\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__38579\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_3\
        );

    \I__7589\ : InMux
    port map (
            O => \N__38574\,
            I => \N__38571\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__38571\,
            I => \phase_controller_inst2.stoper_hc.counter_i_3\
        );

    \I__7587\ : InMux
    port map (
            O => \N__38568\,
            I => \N__38564\
        );

    \I__7586\ : InMux
    port map (
            O => \N__38567\,
            I => \N__38561\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__38564\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_4\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__38561\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_4\
        );

    \I__7583\ : InMux
    port map (
            O => \N__38556\,
            I => \N__38553\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__38553\,
            I => \phase_controller_inst2.stoper_hc.counter_i_4\
        );

    \I__7581\ : InMux
    port map (
            O => \N__38550\,
            I => \N__38546\
        );

    \I__7580\ : InMux
    port map (
            O => \N__38549\,
            I => \N__38543\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__38546\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_5\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__38543\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_5\
        );

    \I__7577\ : CascadeMux
    port map (
            O => \N__38538\,
            I => \N__38535\
        );

    \I__7576\ : InMux
    port map (
            O => \N__38535\,
            I => \N__38532\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__38532\,
            I => \phase_controller_inst2.stoper_hc.counter_i_5\
        );

    \I__7574\ : InMux
    port map (
            O => \N__38529\,
            I => \N__38525\
        );

    \I__7573\ : InMux
    port map (
            O => \N__38528\,
            I => \N__38522\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__38525\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_6\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__38522\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_6\
        );

    \I__7570\ : CascadeMux
    port map (
            O => \N__38517\,
            I => \N__38514\
        );

    \I__7569\ : InMux
    port map (
            O => \N__38514\,
            I => \N__38511\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__38511\,
            I => \N__38508\
        );

    \I__7567\ : Odrv4
    port map (
            O => \N__38508\,
            I => \phase_controller_inst2.stoper_hc.counter_i_6\
        );

    \I__7566\ : InMux
    port map (
            O => \N__38505\,
            I => \N__38501\
        );

    \I__7565\ : InMux
    port map (
            O => \N__38504\,
            I => \N__38498\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__38501\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_7\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__38498\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_7\
        );

    \I__7562\ : CascadeMux
    port map (
            O => \N__38493\,
            I => \N__38490\
        );

    \I__7561\ : InMux
    port map (
            O => \N__38490\,
            I => \N__38487\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__38487\,
            I => \phase_controller_inst2.stoper_hc.counter_i_7\
        );

    \I__7559\ : InMux
    port map (
            O => \N__38484\,
            I => \N__38480\
        );

    \I__7558\ : InMux
    port map (
            O => \N__38483\,
            I => \N__38477\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__38480\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_8\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__38477\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_8\
        );

    \I__7555\ : CascadeMux
    port map (
            O => \N__38472\,
            I => \N__38469\
        );

    \I__7554\ : InMux
    port map (
            O => \N__38469\,
            I => \N__38466\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__38466\,
            I => \phase_controller_inst2.stoper_hc.counter_i_8\
        );

    \I__7552\ : InMux
    port map (
            O => \N__38463\,
            I => \N__38459\
        );

    \I__7551\ : InMux
    port map (
            O => \N__38462\,
            I => \N__38456\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__38459\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_9\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__38456\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_9\
        );

    \I__7548\ : CascadeMux
    port map (
            O => \N__38451\,
            I => \N__38448\
        );

    \I__7547\ : InMux
    port map (
            O => \N__38448\,
            I => \N__38445\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__38445\,
            I => \phase_controller_inst2.stoper_hc.counter_i_9\
        );

    \I__7545\ : InMux
    port map (
            O => \N__38442\,
            I => \N__38438\
        );

    \I__7544\ : InMux
    port map (
            O => \N__38441\,
            I => \N__38435\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__38438\,
            I => \N__38432\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__38435\,
            I => \N__38429\
        );

    \I__7541\ : Odrv12
    port map (
            O => \N__38432\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_19
        );

    \I__7540\ : Odrv12
    port map (
            O => \N__38429\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_19
        );

    \I__7539\ : CEMux
    port map (
            O => \N__38424\,
            I => \N__38420\
        );

    \I__7538\ : CEMux
    port map (
            O => \N__38423\,
            I => \N__38416\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__38420\,
            I => \N__38413\
        );

    \I__7536\ : CEMux
    port map (
            O => \N__38419\,
            I => \N__38410\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__38416\,
            I => \N__38406\
        );

    \I__7534\ : Span4Mux_h
    port map (
            O => \N__38413\,
            I => \N__38401\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__38410\,
            I => \N__38398\
        );

    \I__7532\ : CEMux
    port map (
            O => \N__38409\,
            I => \N__38395\
        );

    \I__7531\ : Span4Mux_v
    port map (
            O => \N__38406\,
            I => \N__38392\
        );

    \I__7530\ : CEMux
    port map (
            O => \N__38405\,
            I => \N__38389\
        );

    \I__7529\ : CEMux
    port map (
            O => \N__38404\,
            I => \N__38386\
        );

    \I__7528\ : Span4Mux_v
    port map (
            O => \N__38401\,
            I => \N__38375\
        );

    \I__7527\ : Span4Mux_v
    port map (
            O => \N__38398\,
            I => \N__38375\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__38395\,
            I => \N__38375\
        );

    \I__7525\ : Span4Mux_v
    port map (
            O => \N__38392\,
            I => \N__38375\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__38389\,
            I => \N__38375\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__38386\,
            I => \N__38371\
        );

    \I__7522\ : Span4Mux_v
    port map (
            O => \N__38375\,
            I => \N__38368\
        );

    \I__7521\ : CEMux
    port map (
            O => \N__38374\,
            I => \N__38365\
        );

    \I__7520\ : Odrv12
    port map (
            O => \N__38371\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__7519\ : Odrv4
    port map (
            O => \N__38368\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__38365\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__7517\ : CascadeMux
    port map (
            O => \N__38358\,
            I => \N__38355\
        );

    \I__7516\ : InMux
    port map (
            O => \N__38355\,
            I => \N__38352\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__38352\,
            I => \N__38349\
        );

    \I__7514\ : Span4Mux_h
    port map (
            O => \N__38349\,
            I => \N__38346\
        );

    \I__7513\ : Odrv4
    port map (
            O => \N__38346\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18\
        );

    \I__7512\ : InMux
    port map (
            O => \N__38343\,
            I => \N__38338\
        );

    \I__7511\ : InMux
    port map (
            O => \N__38342\,
            I => \N__38333\
        );

    \I__7510\ : InMux
    port map (
            O => \N__38341\,
            I => \N__38333\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__38338\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_18\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__38333\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_18\
        );

    \I__7507\ : InMux
    port map (
            O => \N__38328\,
            I => \N__38322\
        );

    \I__7506\ : InMux
    port map (
            O => \N__38327\,
            I => \N__38322\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__38322\,
            I => \N__38319\
        );

    \I__7504\ : Span4Mux_v
    port map (
            O => \N__38319\,
            I => \N__38316\
        );

    \I__7503\ : Odrv4
    port map (
            O => \N__38316\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_18\
        );

    \I__7502\ : CascadeMux
    port map (
            O => \N__38313\,
            I => \N__38309\
        );

    \I__7501\ : InMux
    port map (
            O => \N__38312\,
            I => \N__38304\
        );

    \I__7500\ : InMux
    port map (
            O => \N__38309\,
            I => \N__38304\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__38304\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_19\
        );

    \I__7498\ : CascadeMux
    port map (
            O => \N__38301\,
            I => \N__38296\
        );

    \I__7497\ : InMux
    port map (
            O => \N__38300\,
            I => \N__38293\
        );

    \I__7496\ : InMux
    port map (
            O => \N__38299\,
            I => \N__38288\
        );

    \I__7495\ : InMux
    port map (
            O => \N__38296\,
            I => \N__38288\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__38293\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_19\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__38288\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_19\
        );

    \I__7492\ : InMux
    port map (
            O => \N__38283\,
            I => \N__38280\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__38280\,
            I => \N__38277\
        );

    \I__7490\ : Span4Mux_h
    port map (
            O => \N__38277\,
            I => \N__38274\
        );

    \I__7489\ : Odrv4
    port map (
            O => \N__38274\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt18\
        );

    \I__7488\ : InMux
    port map (
            O => \N__38271\,
            I => \N__38268\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__38268\,
            I => \N__38265\
        );

    \I__7486\ : Span4Mux_s2_v
    port map (
            O => \N__38265\,
            I => \N__38262\
        );

    \I__7485\ : Span4Mux_v
    port map (
            O => \N__38262\,
            I => \N__38257\
        );

    \I__7484\ : InMux
    port map (
            O => \N__38261\,
            I => \N__38252\
        );

    \I__7483\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38252\
        );

    \I__7482\ : Span4Mux_v
    port map (
            O => \N__38257\,
            I => \N__38247\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__38252\,
            I => \N__38247\
        );

    \I__7480\ : Span4Mux_v
    port map (
            O => \N__38247\,
            I => \N__38243\
        );

    \I__7479\ : InMux
    port map (
            O => \N__38246\,
            I => \N__38240\
        );

    \I__7478\ : Odrv4
    port map (
            O => \N__38243\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__38240\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7476\ : IoInMux
    port map (
            O => \N__38235\,
            I => \N__38232\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__38232\,
            I => \N__38229\
        );

    \I__7474\ : Odrv12
    port map (
            O => \N__38229\,
            I => s2_phy_c
        );

    \I__7473\ : IoInMux
    port map (
            O => \N__38226\,
            I => \N__38223\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__38223\,
            I => \current_shift_inst.timer_s1.N_153_i\
        );

    \I__7471\ : CascadeMux
    port map (
            O => \N__38220\,
            I => \N__38216\
        );

    \I__7470\ : InMux
    port map (
            O => \N__38219\,
            I => \N__38209\
        );

    \I__7469\ : InMux
    port map (
            O => \N__38216\,
            I => \N__38206\
        );

    \I__7468\ : InMux
    port map (
            O => \N__38215\,
            I => \N__38203\
        );

    \I__7467\ : InMux
    port map (
            O => \N__38214\,
            I => \N__38200\
        );

    \I__7466\ : InMux
    port map (
            O => \N__38213\,
            I => \N__38197\
        );

    \I__7465\ : CascadeMux
    port map (
            O => \N__38212\,
            I => \N__38194\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__38209\,
            I => \N__38191\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__38206\,
            I => \N__38182\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__38203\,
            I => \N__38182\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__38200\,
            I => \N__38182\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__38197\,
            I => \N__38182\
        );

    \I__7459\ : InMux
    port map (
            O => \N__38194\,
            I => \N__38179\
        );

    \I__7458\ : Span4Mux_h
    port map (
            O => \N__38191\,
            I => \N__38176\
        );

    \I__7457\ : Odrv4
    port map (
            O => \N__38182\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__38179\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__7455\ : Odrv4
    port map (
            O => \N__38176\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__7454\ : CascadeMux
    port map (
            O => \N__38169\,
            I => \N__38166\
        );

    \I__7453\ : InMux
    port map (
            O => \N__38166\,
            I => \N__38162\
        );

    \I__7452\ : InMux
    port map (
            O => \N__38165\,
            I => \N__38159\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__38162\,
            I => \N__38156\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__38159\,
            I => \phase_controller_inst2.stoper_hc.counter\
        );

    \I__7449\ : Odrv4
    port map (
            O => \N__38156\,
            I => \phase_controller_inst2.stoper_hc.counter\
        );

    \I__7448\ : InMux
    port map (
            O => \N__38151\,
            I => \N__38147\
        );

    \I__7447\ : InMux
    port map (
            O => \N__38150\,
            I => \N__38144\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__38147\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_0\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__38144\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_0\
        );

    \I__7444\ : InMux
    port map (
            O => \N__38139\,
            I => \N__38136\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__38136\,
            I => \phase_controller_inst2.stoper_hc.counter_i_0\
        );

    \I__7442\ : InMux
    port map (
            O => \N__38133\,
            I => \N__38129\
        );

    \I__7441\ : InMux
    port map (
            O => \N__38132\,
            I => \N__38126\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__38129\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_1\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__38126\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_1\
        );

    \I__7438\ : InMux
    port map (
            O => \N__38121\,
            I => \N__38118\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__38118\,
            I => \phase_controller_inst2.stoper_hc.counter_i_1\
        );

    \I__7436\ : InMux
    port map (
            O => \N__38115\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__7435\ : InMux
    port map (
            O => \N__38112\,
            I => \bfn_13_26_0_\
        );

    \I__7434\ : InMux
    port map (
            O => \N__38109\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__7433\ : InMux
    port map (
            O => \N__38106\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__7432\ : InMux
    port map (
            O => \N__38103\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__7431\ : InMux
    port map (
            O => \N__38100\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__7430\ : InMux
    port map (
            O => \N__38097\,
            I => \N__38067\
        );

    \I__7429\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38067\
        );

    \I__7428\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38058\
        );

    \I__7427\ : InMux
    port map (
            O => \N__38094\,
            I => \N__38058\
        );

    \I__7426\ : InMux
    port map (
            O => \N__38093\,
            I => \N__38058\
        );

    \I__7425\ : InMux
    port map (
            O => \N__38092\,
            I => \N__38058\
        );

    \I__7424\ : InMux
    port map (
            O => \N__38091\,
            I => \N__38045\
        );

    \I__7423\ : InMux
    port map (
            O => \N__38090\,
            I => \N__38045\
        );

    \I__7422\ : InMux
    port map (
            O => \N__38089\,
            I => \N__38045\
        );

    \I__7421\ : InMux
    port map (
            O => \N__38088\,
            I => \N__38045\
        );

    \I__7420\ : InMux
    port map (
            O => \N__38087\,
            I => \N__38036\
        );

    \I__7419\ : InMux
    port map (
            O => \N__38086\,
            I => \N__38036\
        );

    \I__7418\ : InMux
    port map (
            O => \N__38085\,
            I => \N__38036\
        );

    \I__7417\ : InMux
    port map (
            O => \N__38084\,
            I => \N__38036\
        );

    \I__7416\ : InMux
    port map (
            O => \N__38083\,
            I => \N__38027\
        );

    \I__7415\ : InMux
    port map (
            O => \N__38082\,
            I => \N__38027\
        );

    \I__7414\ : InMux
    port map (
            O => \N__38081\,
            I => \N__38027\
        );

    \I__7413\ : InMux
    port map (
            O => \N__38080\,
            I => \N__38027\
        );

    \I__7412\ : InMux
    port map (
            O => \N__38079\,
            I => \N__38018\
        );

    \I__7411\ : InMux
    port map (
            O => \N__38078\,
            I => \N__38018\
        );

    \I__7410\ : InMux
    port map (
            O => \N__38077\,
            I => \N__38018\
        );

    \I__7409\ : InMux
    port map (
            O => \N__38076\,
            I => \N__38018\
        );

    \I__7408\ : InMux
    port map (
            O => \N__38075\,
            I => \N__38009\
        );

    \I__7407\ : InMux
    port map (
            O => \N__38074\,
            I => \N__38009\
        );

    \I__7406\ : InMux
    port map (
            O => \N__38073\,
            I => \N__38009\
        );

    \I__7405\ : InMux
    port map (
            O => \N__38072\,
            I => \N__38009\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__38067\,
            I => \N__38004\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__38058\,
            I => \N__38004\
        );

    \I__7402\ : InMux
    port map (
            O => \N__38057\,
            I => \N__37995\
        );

    \I__7401\ : InMux
    port map (
            O => \N__38056\,
            I => \N__37995\
        );

    \I__7400\ : InMux
    port map (
            O => \N__38055\,
            I => \N__37995\
        );

    \I__7399\ : InMux
    port map (
            O => \N__38054\,
            I => \N__37995\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__38045\,
            I => \N__37982\
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__38036\,
            I => \N__37982\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__38027\,
            I => \N__37982\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__38018\,
            I => \N__37982\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__38009\,
            I => \N__37982\
        );

    \I__7393\ : Span4Mux_v
    port map (
            O => \N__38004\,
            I => \N__37982\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__37995\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7391\ : Odrv4
    port map (
            O => \N__37982\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7390\ : InMux
    port map (
            O => \N__37977\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__7389\ : CEMux
    port map (
            O => \N__37974\,
            I => \N__37969\
        );

    \I__7388\ : CEMux
    port map (
            O => \N__37973\,
            I => \N__37965\
        );

    \I__7387\ : CEMux
    port map (
            O => \N__37972\,
            I => \N__37962\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__37969\,
            I => \N__37959\
        );

    \I__7385\ : CEMux
    port map (
            O => \N__37968\,
            I => \N__37956\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__37965\,
            I => \N__37951\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__37962\,
            I => \N__37951\
        );

    \I__7382\ : Span4Mux_v
    port map (
            O => \N__37959\,
            I => \N__37946\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__37956\,
            I => \N__37946\
        );

    \I__7380\ : Span4Mux_v
    port map (
            O => \N__37951\,
            I => \N__37943\
        );

    \I__7379\ : Span4Mux_v
    port map (
            O => \N__37946\,
            I => \N__37940\
        );

    \I__7378\ : Span4Mux_h
    port map (
            O => \N__37943\,
            I => \N__37937\
        );

    \I__7377\ : Odrv4
    port map (
            O => \N__37940\,
            I => \delay_measurement_inst.delay_tr_timer.N_158_i\
        );

    \I__7376\ : Odrv4
    port map (
            O => \N__37937\,
            I => \delay_measurement_inst.delay_tr_timer.N_158_i\
        );

    \I__7375\ : InMux
    port map (
            O => \N__37932\,
            I => \N__37929\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__37929\,
            I => \N__37926\
        );

    \I__7373\ : Odrv4
    port map (
            O => \N__37926\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt16\
        );

    \I__7372\ : InMux
    port map (
            O => \N__37923\,
            I => \N__37916\
        );

    \I__7371\ : InMux
    port map (
            O => \N__37922\,
            I => \N__37916\
        );

    \I__7370\ : InMux
    port map (
            O => \N__37921\,
            I => \N__37913\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__37916\,
            I => \N__37910\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__37913\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_17\
        );

    \I__7367\ : Odrv4
    port map (
            O => \N__37910\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_17\
        );

    \I__7366\ : InMux
    port map (
            O => \N__37905\,
            I => \N__37899\
        );

    \I__7365\ : InMux
    port map (
            O => \N__37904\,
            I => \N__37899\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__37899\,
            I => \N__37896\
        );

    \I__7363\ : Span4Mux_v
    port map (
            O => \N__37896\,
            I => \N__37893\
        );

    \I__7362\ : Odrv4
    port map (
            O => \N__37893\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16\
        );

    \I__7361\ : CascadeMux
    port map (
            O => \N__37890\,
            I => \N__37886\
        );

    \I__7360\ : CascadeMux
    port map (
            O => \N__37889\,
            I => \N__37883\
        );

    \I__7359\ : InMux
    port map (
            O => \N__37886\,
            I => \N__37878\
        );

    \I__7358\ : InMux
    port map (
            O => \N__37883\,
            I => \N__37878\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__37878\,
            I => \N__37875\
        );

    \I__7356\ : Span4Mux_v
    port map (
            O => \N__37875\,
            I => \N__37872\
        );

    \I__7355\ : Odrv4
    port map (
            O => \N__37872\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17\
        );

    \I__7354\ : InMux
    port map (
            O => \N__37869\,
            I => \N__37862\
        );

    \I__7353\ : InMux
    port map (
            O => \N__37868\,
            I => \N__37862\
        );

    \I__7352\ : InMux
    port map (
            O => \N__37867\,
            I => \N__37859\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__37862\,
            I => \N__37856\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__37859\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_16\
        );

    \I__7349\ : Odrv4
    port map (
            O => \N__37856\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_16\
        );

    \I__7348\ : CascadeMux
    port map (
            O => \N__37851\,
            I => \N__37848\
        );

    \I__7347\ : InMux
    port map (
            O => \N__37848\,
            I => \N__37845\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__37845\,
            I => \N__37842\
        );

    \I__7345\ : Odrv4
    port map (
            O => \N__37842\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16\
        );

    \I__7344\ : InMux
    port map (
            O => \N__37839\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__7343\ : InMux
    port map (
            O => \N__37836\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__7342\ : InMux
    port map (
            O => \N__37833\,
            I => \bfn_13_25_0_\
        );

    \I__7341\ : InMux
    port map (
            O => \N__37830\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__7340\ : InMux
    port map (
            O => \N__37827\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__7339\ : InMux
    port map (
            O => \N__37824\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__7338\ : InMux
    port map (
            O => \N__37821\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__7337\ : InMux
    port map (
            O => \N__37818\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__7336\ : InMux
    port map (
            O => \N__37815\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__7335\ : InMux
    port map (
            O => \N__37812\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__7334\ : InMux
    port map (
            O => \N__37809\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__7333\ : InMux
    port map (
            O => \N__37806\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__7332\ : InMux
    port map (
            O => \N__37803\,
            I => \bfn_13_24_0_\
        );

    \I__7331\ : InMux
    port map (
            O => \N__37800\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__7330\ : InMux
    port map (
            O => \N__37797\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__7329\ : InMux
    port map (
            O => \N__37794\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__7328\ : InMux
    port map (
            O => \N__37791\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__7327\ : InMux
    port map (
            O => \N__37788\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__7326\ : InMux
    port map (
            O => \N__37785\,
            I => \N__37782\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__37782\,
            I => \N__37779\
        );

    \I__7324\ : Span12Mux_v
    port map (
            O => \N__37779\,
            I => \N__37775\
        );

    \I__7323\ : InMux
    port map (
            O => \N__37778\,
            I => \N__37772\
        );

    \I__7322\ : Odrv12
    port map (
            O => \N__37775\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_26
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__37772\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_26
        );

    \I__7320\ : InMux
    port map (
            O => \N__37767\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25\
        );

    \I__7319\ : InMux
    port map (
            O => \N__37764\,
            I => \N__37761\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__37761\,
            I => \N__37758\
        );

    \I__7317\ : Span12Mux_v
    port map (
            O => \N__37758\,
            I => \N__37754\
        );

    \I__7316\ : InMux
    port map (
            O => \N__37757\,
            I => \N__37751\
        );

    \I__7315\ : Odrv12
    port map (
            O => \N__37754\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_27
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__37751\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_27
        );

    \I__7313\ : InMux
    port map (
            O => \N__37746\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26\
        );

    \I__7312\ : InMux
    port map (
            O => \N__37743\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27\
        );

    \I__7311\ : InMux
    port map (
            O => \N__37740\,
            I => \N__37734\
        );

    \I__7310\ : InMux
    port map (
            O => \N__37739\,
            I => \N__37731\
        );

    \I__7309\ : InMux
    port map (
            O => \N__37738\,
            I => \N__37728\
        );

    \I__7308\ : InMux
    port map (
            O => \N__37737\,
            I => \N__37725\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__37734\,
            I => \N__37720\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__37731\,
            I => \N__37720\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__37728\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__37725\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7303\ : Odrv12
    port map (
            O => \N__37720\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7302\ : InMux
    port map (
            O => \N__37713\,
            I => \bfn_13_23_0_\
        );

    \I__7301\ : InMux
    port map (
            O => \N__37710\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__7300\ : InMux
    port map (
            O => \N__37707\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__7299\ : InMux
    port map (
            O => \N__37704\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__7298\ : InMux
    port map (
            O => \N__37701\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__7297\ : InMux
    port map (
            O => \N__37698\,
            I => \N__37695\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__37695\,
            I => \N__37691\
        );

    \I__7295\ : InMux
    port map (
            O => \N__37694\,
            I => \N__37688\
        );

    \I__7294\ : Odrv12
    port map (
            O => \N__37691\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_18
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__37688\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_18
        );

    \I__7292\ : InMux
    port map (
            O => \N__37683\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17\
        );

    \I__7291\ : InMux
    port map (
            O => \N__37680\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18\
        );

    \I__7290\ : InMux
    port map (
            O => \N__37677\,
            I => \N__37673\
        );

    \I__7289\ : InMux
    port map (
            O => \N__37676\,
            I => \N__37670\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__37673\,
            I => \N__37667\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__37670\,
            I => \N__37664\
        );

    \I__7286\ : Sp12to4
    port map (
            O => \N__37667\,
            I => \N__37661\
        );

    \I__7285\ : Odrv4
    port map (
            O => \N__37664\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_20
        );

    \I__7284\ : Odrv12
    port map (
            O => \N__37661\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_20
        );

    \I__7283\ : InMux
    port map (
            O => \N__37656\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19\
        );

    \I__7282\ : InMux
    port map (
            O => \N__37653\,
            I => \N__37650\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__37650\,
            I => \N__37647\
        );

    \I__7280\ : Span12Mux_v
    port map (
            O => \N__37647\,
            I => \N__37643\
        );

    \I__7279\ : InMux
    port map (
            O => \N__37646\,
            I => \N__37640\
        );

    \I__7278\ : Odrv12
    port map (
            O => \N__37643\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_21
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__37640\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_21
        );

    \I__7276\ : InMux
    port map (
            O => \N__37635\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20\
        );

    \I__7275\ : InMux
    port map (
            O => \N__37632\,
            I => \N__37629\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__37629\,
            I => \N__37626\
        );

    \I__7273\ : Span12Mux_v
    port map (
            O => \N__37626\,
            I => \N__37622\
        );

    \I__7272\ : InMux
    port map (
            O => \N__37625\,
            I => \N__37619\
        );

    \I__7271\ : Odrv12
    port map (
            O => \N__37622\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_22
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__37619\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_22
        );

    \I__7269\ : InMux
    port map (
            O => \N__37614\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21\
        );

    \I__7268\ : InMux
    port map (
            O => \N__37611\,
            I => \N__37608\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__37608\,
            I => \N__37605\
        );

    \I__7266\ : Span12Mux_v
    port map (
            O => \N__37605\,
            I => \N__37601\
        );

    \I__7265\ : InMux
    port map (
            O => \N__37604\,
            I => \N__37598\
        );

    \I__7264\ : Odrv12
    port map (
            O => \N__37601\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_23
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__37598\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_23
        );

    \I__7262\ : InMux
    port map (
            O => \N__37593\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22\
        );

    \I__7261\ : InMux
    port map (
            O => \N__37590\,
            I => \N__37587\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__37587\,
            I => \N__37584\
        );

    \I__7259\ : Sp12to4
    port map (
            O => \N__37584\,
            I => \N__37580\
        );

    \I__7258\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37577\
        );

    \I__7257\ : Odrv12
    port map (
            O => \N__37580\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_24
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__37577\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_24
        );

    \I__7255\ : InMux
    port map (
            O => \N__37572\,
            I => \bfn_13_22_0_\
        );

    \I__7254\ : InMux
    port map (
            O => \N__37569\,
            I => \N__37566\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__37566\,
            I => \N__37563\
        );

    \I__7252\ : Sp12to4
    port map (
            O => \N__37563\,
            I => \N__37559\
        );

    \I__7251\ : InMux
    port map (
            O => \N__37562\,
            I => \N__37556\
        );

    \I__7250\ : Odrv12
    port map (
            O => \N__37559\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_25
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__37556\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_25
        );

    \I__7248\ : InMux
    port map (
            O => \N__37551\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24\
        );

    \I__7247\ : InMux
    port map (
            O => \N__37548\,
            I => \N__37545\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__37545\,
            I => \N__37542\
        );

    \I__7245\ : Span4Mux_v
    port map (
            O => \N__37542\,
            I => \N__37538\
        );

    \I__7244\ : InMux
    port map (
            O => \N__37541\,
            I => \N__37535\
        );

    \I__7243\ : Span4Mux_v
    port map (
            O => \N__37538\,
            I => \N__37530\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__37535\,
            I => \N__37530\
        );

    \I__7241\ : Odrv4
    port map (
            O => \N__37530\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_9
        );

    \I__7240\ : InMux
    port map (
            O => \N__37527\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8\
        );

    \I__7239\ : InMux
    port map (
            O => \N__37524\,
            I => \N__37521\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__37521\,
            I => \N__37518\
        );

    \I__7237\ : Span4Mux_v
    port map (
            O => \N__37518\,
            I => \N__37514\
        );

    \I__7236\ : InMux
    port map (
            O => \N__37517\,
            I => \N__37511\
        );

    \I__7235\ : Odrv4
    port map (
            O => \N__37514\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_10
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__37511\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_10
        );

    \I__7233\ : InMux
    port map (
            O => \N__37506\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9\
        );

    \I__7232\ : InMux
    port map (
            O => \N__37503\,
            I => \N__37500\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__37500\,
            I => \N__37497\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__37497\,
            I => \N__37493\
        );

    \I__7229\ : InMux
    port map (
            O => \N__37496\,
            I => \N__37490\
        );

    \I__7228\ : Odrv4
    port map (
            O => \N__37493\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_11
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__37490\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_11
        );

    \I__7226\ : InMux
    port map (
            O => \N__37485\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10\
        );

    \I__7225\ : InMux
    port map (
            O => \N__37482\,
            I => \N__37479\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__37479\,
            I => \N__37476\
        );

    \I__7223\ : Span4Mux_v
    port map (
            O => \N__37476\,
            I => \N__37472\
        );

    \I__7222\ : InMux
    port map (
            O => \N__37475\,
            I => \N__37469\
        );

    \I__7221\ : Odrv4
    port map (
            O => \N__37472\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_12
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__37469\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_12
        );

    \I__7219\ : InMux
    port map (
            O => \N__37464\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11\
        );

    \I__7218\ : InMux
    port map (
            O => \N__37461\,
            I => \N__37458\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__37458\,
            I => \N__37455\
        );

    \I__7216\ : Span12Mux_v
    port map (
            O => \N__37455\,
            I => \N__37451\
        );

    \I__7215\ : InMux
    port map (
            O => \N__37454\,
            I => \N__37448\
        );

    \I__7214\ : Odrv12
    port map (
            O => \N__37451\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_13
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__37448\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_13
        );

    \I__7212\ : InMux
    port map (
            O => \N__37443\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12\
        );

    \I__7211\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37437\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__37437\,
            I => \N__37434\
        );

    \I__7209\ : Span4Mux_v
    port map (
            O => \N__37434\,
            I => \N__37430\
        );

    \I__7208\ : InMux
    port map (
            O => \N__37433\,
            I => \N__37427\
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__37430\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_14
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__37427\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_14
        );

    \I__7205\ : InMux
    port map (
            O => \N__37422\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13\
        );

    \I__7204\ : InMux
    port map (
            O => \N__37419\,
            I => \N__37416\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__37416\,
            I => \N__37413\
        );

    \I__7202\ : Span12Mux_v
    port map (
            O => \N__37413\,
            I => \N__37409\
        );

    \I__7201\ : InMux
    port map (
            O => \N__37412\,
            I => \N__37406\
        );

    \I__7200\ : Odrv12
    port map (
            O => \N__37409\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_15
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__37406\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_15
        );

    \I__7198\ : InMux
    port map (
            O => \N__37401\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14\
        );

    \I__7197\ : InMux
    port map (
            O => \N__37398\,
            I => \N__37395\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__37395\,
            I => \N__37392\
        );

    \I__7195\ : Span12Mux_v
    port map (
            O => \N__37392\,
            I => \N__37388\
        );

    \I__7194\ : InMux
    port map (
            O => \N__37391\,
            I => \N__37385\
        );

    \I__7193\ : Odrv12
    port map (
            O => \N__37388\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_16
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__37385\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_16
        );

    \I__7191\ : InMux
    port map (
            O => \N__37380\,
            I => \bfn_13_21_0_\
        );

    \I__7190\ : InMux
    port map (
            O => \N__37377\,
            I => \N__37374\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__37374\,
            I => \N__37370\
        );

    \I__7188\ : InMux
    port map (
            O => \N__37373\,
            I => \N__37367\
        );

    \I__7187\ : Sp12to4
    port map (
            O => \N__37370\,
            I => \N__37364\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__37367\,
            I => \N__37361\
        );

    \I__7185\ : Odrv12
    port map (
            O => \N__37364\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_17
        );

    \I__7184\ : Odrv4
    port map (
            O => \N__37361\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_17
        );

    \I__7183\ : InMux
    port map (
            O => \N__37356\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16\
        );

    \I__7182\ : InMux
    port map (
            O => \N__37353\,
            I => \N__37349\
        );

    \I__7181\ : InMux
    port map (
            O => \N__37352\,
            I => \N__37346\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__37349\,
            I => \N__37343\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__37346\,
            I => \N__37340\
        );

    \I__7178\ : Sp12to4
    port map (
            O => \N__37343\,
            I => \N__37337\
        );

    \I__7177\ : Span4Mux_v
    port map (
            O => \N__37340\,
            I => \N__37334\
        );

    \I__7176\ : Span12Mux_s7_v
    port map (
            O => \N__37337\,
            I => \N__37331\
        );

    \I__7175\ : Odrv4
    port map (
            O => \N__37334\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_1
        );

    \I__7174\ : Odrv12
    port map (
            O => \N__37331\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_1
        );

    \I__7173\ : InMux
    port map (
            O => \N__37326\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0\
        );

    \I__7172\ : InMux
    port map (
            O => \N__37323\,
            I => \N__37320\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__37320\,
            I => \N__37316\
        );

    \I__7170\ : InMux
    port map (
            O => \N__37319\,
            I => \N__37313\
        );

    \I__7169\ : Span12Mux_h
    port map (
            O => \N__37316\,
            I => \N__37310\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__37313\,
            I => \N__37307\
        );

    \I__7167\ : Span12Mux_v
    port map (
            O => \N__37310\,
            I => \N__37304\
        );

    \I__7166\ : Span4Mux_v
    port map (
            O => \N__37307\,
            I => \N__37301\
        );

    \I__7165\ : Odrv12
    port map (
            O => \N__37304\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_2
        );

    \I__7164\ : Odrv4
    port map (
            O => \N__37301\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_2
        );

    \I__7163\ : InMux
    port map (
            O => \N__37296\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1\
        );

    \I__7162\ : InMux
    port map (
            O => \N__37293\,
            I => \N__37290\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__37290\,
            I => \N__37286\
        );

    \I__7160\ : InMux
    port map (
            O => \N__37289\,
            I => \N__37283\
        );

    \I__7159\ : Sp12to4
    port map (
            O => \N__37286\,
            I => \N__37280\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__37283\,
            I => \N__37277\
        );

    \I__7157\ : Span12Mux_v
    port map (
            O => \N__37280\,
            I => \N__37274\
        );

    \I__7156\ : Span4Mux_v
    port map (
            O => \N__37277\,
            I => \N__37271\
        );

    \I__7155\ : Odrv12
    port map (
            O => \N__37274\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_3
        );

    \I__7154\ : Odrv4
    port map (
            O => \N__37271\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_3
        );

    \I__7153\ : InMux
    port map (
            O => \N__37266\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2\
        );

    \I__7152\ : InMux
    port map (
            O => \N__37263\,
            I => \N__37259\
        );

    \I__7151\ : InMux
    port map (
            O => \N__37262\,
            I => \N__37256\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__37259\,
            I => \N__37253\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__37256\,
            I => \N__37250\
        );

    \I__7148\ : Span4Mux_h
    port map (
            O => \N__37253\,
            I => \N__37247\
        );

    \I__7147\ : Span4Mux_v
    port map (
            O => \N__37250\,
            I => \N__37244\
        );

    \I__7146\ : Span4Mux_v
    port map (
            O => \N__37247\,
            I => \N__37241\
        );

    \I__7145\ : Odrv4
    port map (
            O => \N__37244\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_4
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__37241\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_4
        );

    \I__7143\ : InMux
    port map (
            O => \N__37236\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3\
        );

    \I__7142\ : InMux
    port map (
            O => \N__37233\,
            I => \N__37230\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__37230\,
            I => \N__37226\
        );

    \I__7140\ : InMux
    port map (
            O => \N__37229\,
            I => \N__37223\
        );

    \I__7139\ : Span12Mux_s6_v
    port map (
            O => \N__37226\,
            I => \N__37220\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__37223\,
            I => \N__37217\
        );

    \I__7137\ : Span12Mux_v
    port map (
            O => \N__37220\,
            I => \N__37214\
        );

    \I__7136\ : Span4Mux_v
    port map (
            O => \N__37217\,
            I => \N__37211\
        );

    \I__7135\ : Odrv12
    port map (
            O => \N__37214\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_5
        );

    \I__7134\ : Odrv4
    port map (
            O => \N__37211\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_5
        );

    \I__7133\ : InMux
    port map (
            O => \N__37206\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4\
        );

    \I__7132\ : InMux
    port map (
            O => \N__37203\,
            I => \N__37199\
        );

    \I__7131\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37196\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__37199\,
            I => \N__37193\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__37196\,
            I => \N__37190\
        );

    \I__7128\ : Span4Mux_v
    port map (
            O => \N__37193\,
            I => \N__37187\
        );

    \I__7127\ : Span4Mux_v
    port map (
            O => \N__37190\,
            I => \N__37184\
        );

    \I__7126\ : Odrv4
    port map (
            O => \N__37187\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_6
        );

    \I__7125\ : Odrv4
    port map (
            O => \N__37184\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_6
        );

    \I__7124\ : InMux
    port map (
            O => \N__37179\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5\
        );

    \I__7123\ : InMux
    port map (
            O => \N__37176\,
            I => \N__37173\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__37173\,
            I => \N__37169\
        );

    \I__7121\ : InMux
    port map (
            O => \N__37172\,
            I => \N__37166\
        );

    \I__7120\ : Span4Mux_v
    port map (
            O => \N__37169\,
            I => \N__37163\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__37166\,
            I => \N__37160\
        );

    \I__7118\ : Odrv4
    port map (
            O => \N__37163\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_7
        );

    \I__7117\ : Odrv4
    port map (
            O => \N__37160\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_7
        );

    \I__7116\ : InMux
    port map (
            O => \N__37155\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6\
        );

    \I__7115\ : InMux
    port map (
            O => \N__37152\,
            I => \N__37149\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__37149\,
            I => \N__37145\
        );

    \I__7113\ : InMux
    port map (
            O => \N__37148\,
            I => \N__37142\
        );

    \I__7112\ : Sp12to4
    port map (
            O => \N__37145\,
            I => \N__37139\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__37142\,
            I => \N__37136\
        );

    \I__7110\ : Span12Mux_v
    port map (
            O => \N__37139\,
            I => \N__37133\
        );

    \I__7109\ : Span4Mux_v
    port map (
            O => \N__37136\,
            I => \N__37130\
        );

    \I__7108\ : Odrv12
    port map (
            O => \N__37133\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_8
        );

    \I__7107\ : Odrv4
    port map (
            O => \N__37130\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_8
        );

    \I__7106\ : InMux
    port map (
            O => \N__37125\,
            I => \bfn_13_20_0_\
        );

    \I__7105\ : InMux
    port map (
            O => \N__37122\,
            I => \N__37119\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__37119\,
            I => \N__37116\
        );

    \I__7103\ : Span4Mux_v
    port map (
            O => \N__37116\,
            I => \N__37113\
        );

    \I__7102\ : Span4Mux_h
    port map (
            O => \N__37113\,
            I => \N__37110\
        );

    \I__7101\ : Odrv4
    port map (
            O => \N__37110\,
            I => \phase_controller_inst1.stoper_tr.un4_start_0\
        );

    \I__7100\ : CascadeMux
    port map (
            O => \N__37107\,
            I => \N__37103\
        );

    \I__7099\ : InMux
    port map (
            O => \N__37106\,
            I => \N__37095\
        );

    \I__7098\ : InMux
    port map (
            O => \N__37103\,
            I => \N__37095\
        );

    \I__7097\ : InMux
    port map (
            O => \N__37102\,
            I => \N__37095\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__37095\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__7095\ : InMux
    port map (
            O => \N__37092\,
            I => \N__37086\
        );

    \I__7094\ : InMux
    port map (
            O => \N__37091\,
            I => \N__37086\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__37086\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__7092\ : CascadeMux
    port map (
            O => \N__37083\,
            I => \N__37079\
        );

    \I__7091\ : InMux
    port map (
            O => \N__37082\,
            I => \N__37076\
        );

    \I__7090\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37073\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__37076\,
            I => \N__37067\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__37073\,
            I => \N__37067\
        );

    \I__7087\ : InMux
    port map (
            O => \N__37072\,
            I => \N__37064\
        );

    \I__7086\ : Span4Mux_v
    port map (
            O => \N__37067\,
            I => \N__37059\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__37064\,
            I => \N__37059\
        );

    \I__7084\ : Span4Mux_h
    port map (
            O => \N__37059\,
            I => \N__37056\
        );

    \I__7083\ : Sp12to4
    port map (
            O => \N__37056\,
            I => \N__37053\
        );

    \I__7082\ : Span12Mux_v
    port map (
            O => \N__37053\,
            I => \N__37050\
        );

    \I__7081\ : Odrv12
    port map (
            O => \N__37050\,
            I => il_min_comp1_c
        );

    \I__7080\ : InMux
    port map (
            O => \N__37047\,
            I => \N__37044\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__37044\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa\
        );

    \I__7078\ : InMux
    port map (
            O => \N__37041\,
            I => \N__37037\
        );

    \I__7077\ : InMux
    port map (
            O => \N__37040\,
            I => \N__37033\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__37037\,
            I => \N__37028\
        );

    \I__7075\ : InMux
    port map (
            O => \N__37036\,
            I => \N__37025\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__37033\,
            I => \N__37022\
        );

    \I__7073\ : InMux
    port map (
            O => \N__37032\,
            I => \N__37017\
        );

    \I__7072\ : InMux
    port map (
            O => \N__37031\,
            I => \N__37017\
        );

    \I__7071\ : Span4Mux_v
    port map (
            O => \N__37028\,
            I => \N__37014\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__37025\,
            I => \N__37010\
        );

    \I__7069\ : Span4Mux_h
    port map (
            O => \N__37022\,
            I => \N__37007\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__37017\,
            I => \N__37002\
        );

    \I__7067\ : Span4Mux_h
    port map (
            O => \N__37014\,
            I => \N__37002\
        );

    \I__7066\ : InMux
    port map (
            O => \N__37013\,
            I => \N__36999\
        );

    \I__7065\ : Span4Mux_h
    port map (
            O => \N__37010\,
            I => \N__36996\
        );

    \I__7064\ : Span4Mux_v
    port map (
            O => \N__37007\,
            I => \N__36993\
        );

    \I__7063\ : Sp12to4
    port map (
            O => \N__37002\,
            I => \N__36990\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__36999\,
            I => \N__36985\
        );

    \I__7061\ : Span4Mux_v
    port map (
            O => \N__36996\,
            I => \N__36985\
        );

    \I__7060\ : Odrv4
    port map (
            O => \N__36993\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__7059\ : Odrv12
    port map (
            O => \N__36990\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__7058\ : Odrv4
    port map (
            O => \N__36985\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__7057\ : CascadeMux
    port map (
            O => \N__36978\,
            I => \N__36975\
        );

    \I__7056\ : InMux
    port map (
            O => \N__36975\,
            I => \N__36971\
        );

    \I__7055\ : InMux
    port map (
            O => \N__36974\,
            I => \N__36967\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__36971\,
            I => \N__36963\
        );

    \I__7053\ : InMux
    port map (
            O => \N__36970\,
            I => \N__36960\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__36967\,
            I => \N__36956\
        );

    \I__7051\ : InMux
    port map (
            O => \N__36966\,
            I => \N__36953\
        );

    \I__7050\ : Span4Mux_h
    port map (
            O => \N__36963\,
            I => \N__36950\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__36960\,
            I => \N__36946\
        );

    \I__7048\ : InMux
    port map (
            O => \N__36959\,
            I => \N__36943\
        );

    \I__7047\ : Span4Mux_h
    port map (
            O => \N__36956\,
            I => \N__36940\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__36953\,
            I => \N__36937\
        );

    \I__7045\ : Span4Mux_v
    port map (
            O => \N__36950\,
            I => \N__36934\
        );

    \I__7044\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36931\
        );

    \I__7043\ : Span12Mux_v
    port map (
            O => \N__36946\,
            I => \N__36928\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__36943\,
            I => \N__36921\
        );

    \I__7041\ : Span4Mux_v
    port map (
            O => \N__36940\,
            I => \N__36921\
        );

    \I__7040\ : Span4Mux_s3_v
    port map (
            O => \N__36937\,
            I => \N__36921\
        );

    \I__7039\ : Odrv4
    port map (
            O => \N__36934\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__36931\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__7037\ : Odrv12
    port map (
            O => \N__36928\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__7036\ : Odrv4
    port map (
            O => \N__36921\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__7035\ : InMux
    port map (
            O => \N__36912\,
            I => \N__36906\
        );

    \I__7034\ : InMux
    port map (
            O => \N__36911\,
            I => \N__36906\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__36906\,
            I => \N__36903\
        );

    \I__7032\ : Span4Mux_h
    port map (
            O => \N__36903\,
            I => \N__36900\
        );

    \I__7031\ : Span4Mux_v
    port map (
            O => \N__36900\,
            I => \N__36897\
        );

    \I__7030\ : Span4Mux_v
    port map (
            O => \N__36897\,
            I => \N__36893\
        );

    \I__7029\ : InMux
    port map (
            O => \N__36896\,
            I => \N__36890\
        );

    \I__7028\ : Odrv4
    port map (
            O => \N__36893\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__36890\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__7026\ : InMux
    port map (
            O => \N__36885\,
            I => \N__36882\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__36882\,
            I => \N__36878\
        );

    \I__7024\ : CascadeMux
    port map (
            O => \N__36881\,
            I => \N__36874\
        );

    \I__7023\ : Span4Mux_h
    port map (
            O => \N__36878\,
            I => \N__36871\
        );

    \I__7022\ : InMux
    port map (
            O => \N__36877\,
            I => \N__36866\
        );

    \I__7021\ : InMux
    port map (
            O => \N__36874\,
            I => \N__36866\
        );

    \I__7020\ : Span4Mux_v
    port map (
            O => \N__36871\,
            I => \N__36863\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__36866\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__7018\ : Odrv4
    port map (
            O => \N__36863\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__7017\ : CascadeMux
    port map (
            O => \N__36858\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\
        );

    \I__7016\ : InMux
    port map (
            O => \N__36855\,
            I => \N__36852\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__36852\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\
        );

    \I__7014\ : CascadeMux
    port map (
            O => \N__36849\,
            I => \N__36846\
        );

    \I__7013\ : InMux
    port map (
            O => \N__36846\,
            I => \N__36840\
        );

    \I__7012\ : InMux
    port map (
            O => \N__36845\,
            I => \N__36835\
        );

    \I__7011\ : InMux
    port map (
            O => \N__36844\,
            I => \N__36835\
        );

    \I__7010\ : InMux
    port map (
            O => \N__36843\,
            I => \N__36832\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__36840\,
            I => \N__36829\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__36835\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__36832\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7006\ : Odrv4
    port map (
            O => \N__36829\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7005\ : InMux
    port map (
            O => \N__36822\,
            I => \N__36818\
        );

    \I__7004\ : InMux
    port map (
            O => \N__36821\,
            I => \N__36814\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__36818\,
            I => \N__36811\
        );

    \I__7002\ : InMux
    port map (
            O => \N__36817\,
            I => \N__36808\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__36814\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__36811\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__36808\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__6998\ : InMux
    port map (
            O => \N__36801\,
            I => \N__36798\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__36798\,
            I => \phase_controller_inst1.stoper_tr.measured_delay_tr_i_31\
        );

    \I__6996\ : InMux
    port map (
            O => \N__36795\,
            I => \N__36791\
        );

    \I__6995\ : InMux
    port map (
            O => \N__36794\,
            I => \N__36788\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__36791\,
            I => \N__36784\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__36788\,
            I => \N__36780\
        );

    \I__6992\ : InMux
    port map (
            O => \N__36787\,
            I => \N__36777\
        );

    \I__6991\ : Span4Mux_h
    port map (
            O => \N__36784\,
            I => \N__36774\
        );

    \I__6990\ : InMux
    port map (
            O => \N__36783\,
            I => \N__36771\
        );

    \I__6989\ : Span4Mux_v
    port map (
            O => \N__36780\,
            I => \N__36768\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__36777\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6987\ : Odrv4
    port map (
            O => \N__36774\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__36771\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6985\ : Odrv4
    port map (
            O => \N__36768\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6984\ : InMux
    port map (
            O => \N__36759\,
            I => \N__36755\
        );

    \I__6983\ : CascadeMux
    port map (
            O => \N__36758\,
            I => \N__36750\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__36755\,
            I => \N__36747\
        );

    \I__6981\ : InMux
    port map (
            O => \N__36754\,
            I => \N__36744\
        );

    \I__6980\ : InMux
    port map (
            O => \N__36753\,
            I => \N__36739\
        );

    \I__6979\ : InMux
    port map (
            O => \N__36750\,
            I => \N__36739\
        );

    \I__6978\ : Span4Mux_v
    port map (
            O => \N__36747\,
            I => \N__36736\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__36744\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6976\ : LocalMux
    port map (
            O => \N__36739\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6975\ : Odrv4
    port map (
            O => \N__36736\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6974\ : InMux
    port map (
            O => \N__36729\,
            I => \N__36725\
        );

    \I__6973\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36722\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__36725\,
            I => \N__36719\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__36722\,
            I => \N__36716\
        );

    \I__6970\ : Span12Mux_v
    port map (
            O => \N__36719\,
            I => \N__36713\
        );

    \I__6969\ : Odrv12
    port map (
            O => \N__36716\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__6968\ : Odrv12
    port map (
            O => \N__36713\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__6967\ : CascadeMux
    port map (
            O => \N__36708\,
            I => \N__36704\
        );

    \I__6966\ : InMux
    port map (
            O => \N__36707\,
            I => \N__36701\
        );

    \I__6965\ : InMux
    port map (
            O => \N__36704\,
            I => \N__36698\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__36701\,
            I => \N__36694\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__36698\,
            I => \N__36691\
        );

    \I__6962\ : CascadeMux
    port map (
            O => \N__36697\,
            I => \N__36688\
        );

    \I__6961\ : Span4Mux_v
    port map (
            O => \N__36694\,
            I => \N__36685\
        );

    \I__6960\ : Span4Mux_v
    port map (
            O => \N__36691\,
            I => \N__36682\
        );

    \I__6959\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36678\
        );

    \I__6958\ : Sp12to4
    port map (
            O => \N__36685\,
            I => \N__36673\
        );

    \I__6957\ : Sp12to4
    port map (
            O => \N__36682\,
            I => \N__36673\
        );

    \I__6956\ : InMux
    port map (
            O => \N__36681\,
            I => \N__36670\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__36678\,
            I => \N__36667\
        );

    \I__6954\ : Span12Mux_h
    port map (
            O => \N__36673\,
            I => \N__36664\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__36670\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__6952\ : Odrv12
    port map (
            O => \N__36667\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__6951\ : Odrv12
    port map (
            O => \N__36664\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__6950\ : InMux
    port map (
            O => \N__36657\,
            I => \N__36654\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__36654\,
            I => \N__36650\
        );

    \I__6948\ : InMux
    port map (
            O => \N__36653\,
            I => \N__36647\
        );

    \I__6947\ : Span4Mux_h
    port map (
            O => \N__36650\,
            I => \N__36641\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__36647\,
            I => \N__36641\
        );

    \I__6945\ : InMux
    port map (
            O => \N__36646\,
            I => \N__36638\
        );

    \I__6944\ : Span4Mux_v
    port map (
            O => \N__36641\,
            I => \N__36635\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__36638\,
            I => \N__36632\
        );

    \I__6942\ : Span4Mux_v
    port map (
            O => \N__36635\,
            I => \N__36629\
        );

    \I__6941\ : Span4Mux_v
    port map (
            O => \N__36632\,
            I => \N__36626\
        );

    \I__6940\ : Sp12to4
    port map (
            O => \N__36629\,
            I => \N__36623\
        );

    \I__6939\ : Span4Mux_h
    port map (
            O => \N__36626\,
            I => \N__36620\
        );

    \I__6938\ : Span12Mux_h
    port map (
            O => \N__36623\,
            I => \N__36615\
        );

    \I__6937\ : Sp12to4
    port map (
            O => \N__36620\,
            I => \N__36615\
        );

    \I__6936\ : Odrv12
    port map (
            O => \N__36615\,
            I => il_max_comp1_c
        );

    \I__6935\ : InMux
    port map (
            O => \N__36612\,
            I => \N__36608\
        );

    \I__6934\ : InMux
    port map (
            O => \N__36611\,
            I => \N__36605\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__36608\,
            I => \N__36601\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__36605\,
            I => \N__36598\
        );

    \I__6931\ : InMux
    port map (
            O => \N__36604\,
            I => \N__36595\
        );

    \I__6930\ : Span4Mux_s3_v
    port map (
            O => \N__36601\,
            I => \N__36590\
        );

    \I__6929\ : Span4Mux_s3_v
    port map (
            O => \N__36598\,
            I => \N__36590\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__36595\,
            I => \N__36585\
        );

    \I__6927\ : Span4Mux_h
    port map (
            O => \N__36590\,
            I => \N__36582\
        );

    \I__6926\ : InMux
    port map (
            O => \N__36589\,
            I => \N__36577\
        );

    \I__6925\ : InMux
    port map (
            O => \N__36588\,
            I => \N__36577\
        );

    \I__6924\ : Span4Mux_v
    port map (
            O => \N__36585\,
            I => \N__36574\
        );

    \I__6923\ : Sp12to4
    port map (
            O => \N__36582\,
            I => \N__36571\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__36577\,
            I => \N__36568\
        );

    \I__6921\ : Span4Mux_h
    port map (
            O => \N__36574\,
            I => \N__36562\
        );

    \I__6920\ : Span12Mux_s11_v
    port map (
            O => \N__36571\,
            I => \N__36557\
        );

    \I__6919\ : Sp12to4
    port map (
            O => \N__36568\,
            I => \N__36557\
        );

    \I__6918\ : InMux
    port map (
            O => \N__36567\,
            I => \N__36550\
        );

    \I__6917\ : InMux
    port map (
            O => \N__36566\,
            I => \N__36550\
        );

    \I__6916\ : InMux
    port map (
            O => \N__36565\,
            I => \N__36550\
        );

    \I__6915\ : Sp12to4
    port map (
            O => \N__36562\,
            I => \N__36547\
        );

    \I__6914\ : Span12Mux_v
    port map (
            O => \N__36557\,
            I => \N__36542\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__36550\,
            I => \N__36542\
        );

    \I__6912\ : Span12Mux_v
    port map (
            O => \N__36547\,
            I => \N__36537\
        );

    \I__6911\ : Span12Mux_h
    port map (
            O => \N__36542\,
            I => \N__36537\
        );

    \I__6910\ : Odrv12
    port map (
            O => \N__36537\,
            I => start_stop_c
        );

    \I__6909\ : InMux
    port map (
            O => \N__36534\,
            I => \N__36531\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__36531\,
            I => \N__36526\
        );

    \I__6907\ : InMux
    port map (
            O => \N__36530\,
            I => \N__36521\
        );

    \I__6906\ : InMux
    port map (
            O => \N__36529\,
            I => \N__36521\
        );

    \I__6905\ : Odrv12
    port map (
            O => \N__36526\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__36521\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__6903\ : CascadeMux
    port map (
            O => \N__36516\,
            I => \phase_controller_inst1.state_ns_0_0_1_cascade_\
        );

    \I__6902\ : InMux
    port map (
            O => \N__36513\,
            I => \N__36509\
        );

    \I__6901\ : CascadeMux
    port map (
            O => \N__36512\,
            I => \N__36506\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__36509\,
            I => \N__36502\
        );

    \I__6899\ : InMux
    port map (
            O => \N__36506\,
            I => \N__36497\
        );

    \I__6898\ : InMux
    port map (
            O => \N__36505\,
            I => \N__36497\
        );

    \I__6897\ : Span12Mux_h
    port map (
            O => \N__36502\,
            I => \N__36494\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__36497\,
            I => \phase_controller_inst1.start_flagZ0\
        );

    \I__6895\ : Odrv12
    port map (
            O => \N__36494\,
            I => \phase_controller_inst1.start_flagZ0\
        );

    \I__6894\ : InMux
    port map (
            O => \N__36489\,
            I => \N__36486\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__36486\,
            I => \N__36483\
        );

    \I__6892\ : Span4Mux_h
    port map (
            O => \N__36483\,
            I => \N__36480\
        );

    \I__6891\ : Odrv4
    port map (
            O => \N__36480\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_15\
        );

    \I__6890\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36473\
        );

    \I__6889\ : InMux
    port map (
            O => \N__36476\,
            I => \N__36470\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__36473\,
            I => \N__36467\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__36470\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27\
        );

    \I__6886\ : Odrv4
    port map (
            O => \N__36467\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27\
        );

    \I__6885\ : InMux
    port map (
            O => \N__36462\,
            I => \N__36456\
        );

    \I__6884\ : InMux
    port map (
            O => \N__36461\,
            I => \N__36456\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__36456\,
            I => \N__36453\
        );

    \I__6882\ : Span4Mux_h
    port map (
            O => \N__36453\,
            I => \N__36450\
        );

    \I__6881\ : Odrv4
    port map (
            O => \N__36450\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_20\
        );

    \I__6880\ : CascadeMux
    port map (
            O => \N__36447\,
            I => \N__36443\
        );

    \I__6879\ : CascadeMux
    port map (
            O => \N__36446\,
            I => \N__36440\
        );

    \I__6878\ : InMux
    port map (
            O => \N__36443\,
            I => \N__36435\
        );

    \I__6877\ : InMux
    port map (
            O => \N__36440\,
            I => \N__36435\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__36435\,
            I => \N__36432\
        );

    \I__6875\ : Span4Mux_h
    port map (
            O => \N__36432\,
            I => \N__36429\
        );

    \I__6874\ : Odrv4
    port map (
            O => \N__36429\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_23\
        );

    \I__6873\ : InMux
    port map (
            O => \N__36426\,
            I => \N__36423\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__36423\,
            I => \N__36420\
        );

    \I__6871\ : Span4Mux_v
    port map (
            O => \N__36420\,
            I => \N__36417\
        );

    \I__6870\ : Span4Mux_v
    port map (
            O => \N__36417\,
            I => \N__36414\
        );

    \I__6869\ : Odrv4
    port map (
            O => \N__36414\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_7\
        );

    \I__6868\ : CascadeMux
    port map (
            O => \N__36411\,
            I => \N__36408\
        );

    \I__6867\ : InMux
    port map (
            O => \N__36408\,
            I => \N__36402\
        );

    \I__6866\ : InMux
    port map (
            O => \N__36407\,
            I => \N__36402\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__36402\,
            I => \N__36399\
        );

    \I__6864\ : Span4Mux_h
    port map (
            O => \N__36399\,
            I => \N__36396\
        );

    \I__6863\ : Odrv4
    port map (
            O => \N__36396\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_18\
        );

    \I__6862\ : InMux
    port map (
            O => \N__36393\,
            I => \N__36387\
        );

    \I__6861\ : InMux
    port map (
            O => \N__36392\,
            I => \N__36387\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__36387\,
            I => \N__36384\
        );

    \I__6859\ : Span4Mux_h
    port map (
            O => \N__36384\,
            I => \N__36381\
        );

    \I__6858\ : Odrv4
    port map (
            O => \N__36381\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_16\
        );

    \I__6857\ : CascadeMux
    port map (
            O => \N__36378\,
            I => \N__36374\
        );

    \I__6856\ : InMux
    port map (
            O => \N__36377\,
            I => \N__36369\
        );

    \I__6855\ : InMux
    port map (
            O => \N__36374\,
            I => \N__36369\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__36369\,
            I => \N__36366\
        );

    \I__6853\ : Span4Mux_h
    port map (
            O => \N__36366\,
            I => \N__36363\
        );

    \I__6852\ : Odrv4
    port map (
            O => \N__36363\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_19\
        );

    \I__6851\ : CascadeMux
    port map (
            O => \N__36360\,
            I => \N__36356\
        );

    \I__6850\ : CascadeMux
    port map (
            O => \N__36359\,
            I => \N__36353\
        );

    \I__6849\ : InMux
    port map (
            O => \N__36356\,
            I => \N__36348\
        );

    \I__6848\ : InMux
    port map (
            O => \N__36353\,
            I => \N__36348\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__36348\,
            I => \N__36345\
        );

    \I__6846\ : Span4Mux_v
    port map (
            O => \N__36345\,
            I => \N__36342\
        );

    \I__6845\ : Odrv4
    port map (
            O => \N__36342\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_21\
        );

    \I__6844\ : CEMux
    port map (
            O => \N__36339\,
            I => \N__36336\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__36336\,
            I => \N__36329\
        );

    \I__6842\ : CEMux
    port map (
            O => \N__36335\,
            I => \N__36326\
        );

    \I__6841\ : CEMux
    port map (
            O => \N__36334\,
            I => \N__36321\
        );

    \I__6840\ : CEMux
    port map (
            O => \N__36333\,
            I => \N__36318\
        );

    \I__6839\ : CEMux
    port map (
            O => \N__36332\,
            I => \N__36315\
        );

    \I__6838\ : Span4Mux_h
    port map (
            O => \N__36329\,
            I => \N__36309\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__36326\,
            I => \N__36309\
        );

    \I__6836\ : CEMux
    port map (
            O => \N__36325\,
            I => \N__36306\
        );

    \I__6835\ : CEMux
    port map (
            O => \N__36324\,
            I => \N__36303\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__36321\,
            I => \N__36298\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__36318\,
            I => \N__36298\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__36315\,
            I => \N__36295\
        );

    \I__6831\ : CEMux
    port map (
            O => \N__36314\,
            I => \N__36292\
        );

    \I__6830\ : Span4Mux_v
    port map (
            O => \N__36309\,
            I => \N__36289\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__36306\,
            I => \N__36286\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__36303\,
            I => \N__36283\
        );

    \I__6827\ : Span4Mux_v
    port map (
            O => \N__36298\,
            I => \N__36276\
        );

    \I__6826\ : Span4Mux_v
    port map (
            O => \N__36295\,
            I => \N__36276\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__36292\,
            I => \N__36276\
        );

    \I__6824\ : Span4Mux_h
    port map (
            O => \N__36289\,
            I => \N__36271\
        );

    \I__6823\ : Span4Mux_v
    port map (
            O => \N__36286\,
            I => \N__36271\
        );

    \I__6822\ : Span4Mux_v
    port map (
            O => \N__36283\,
            I => \N__36266\
        );

    \I__6821\ : Span4Mux_v
    port map (
            O => \N__36276\,
            I => \N__36266\
        );

    \I__6820\ : Odrv4
    port map (
            O => \N__36271\,
            I => \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__6819\ : Odrv4
    port map (
            O => \N__36266\,
            I => \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__6818\ : InMux
    port map (
            O => \N__36261\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_25\
        );

    \I__6817\ : InMux
    port map (
            O => \N__36258\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_26\
        );

    \I__6816\ : InMux
    port map (
            O => \N__36255\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_27\
        );

    \I__6815\ : InMux
    port map (
            O => \N__36252\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_28\
        );

    \I__6814\ : InMux
    port map (
            O => \N__36249\,
            I => \N__36244\
        );

    \I__6813\ : InMux
    port map (
            O => \N__36248\,
            I => \N__36239\
        );

    \I__6812\ : InMux
    port map (
            O => \N__36247\,
            I => \N__36239\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__36244\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_30\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__36239\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_30\
        );

    \I__6809\ : InMux
    port map (
            O => \N__36234\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_29\
        );

    \I__6808\ : InMux
    port map (
            O => \N__36231\,
            I => \N__36214\
        );

    \I__6807\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36214\
        );

    \I__6806\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36214\
        );

    \I__6805\ : InMux
    port map (
            O => \N__36228\,
            I => \N__36184\
        );

    \I__6804\ : InMux
    port map (
            O => \N__36227\,
            I => \N__36184\
        );

    \I__6803\ : InMux
    port map (
            O => \N__36226\,
            I => \N__36184\
        );

    \I__6802\ : InMux
    port map (
            O => \N__36225\,
            I => \N__36184\
        );

    \I__6801\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36175\
        );

    \I__6800\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36175\
        );

    \I__6799\ : InMux
    port map (
            O => \N__36222\,
            I => \N__36175\
        );

    \I__6798\ : InMux
    port map (
            O => \N__36221\,
            I => \N__36175\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__36214\,
            I => \N__36172\
        );

    \I__6796\ : InMux
    port map (
            O => \N__36213\,
            I => \N__36163\
        );

    \I__6795\ : InMux
    port map (
            O => \N__36212\,
            I => \N__36163\
        );

    \I__6794\ : InMux
    port map (
            O => \N__36211\,
            I => \N__36163\
        );

    \I__6793\ : InMux
    port map (
            O => \N__36210\,
            I => \N__36163\
        );

    \I__6792\ : InMux
    port map (
            O => \N__36209\,
            I => \N__36154\
        );

    \I__6791\ : InMux
    port map (
            O => \N__36208\,
            I => \N__36154\
        );

    \I__6790\ : InMux
    port map (
            O => \N__36207\,
            I => \N__36154\
        );

    \I__6789\ : InMux
    port map (
            O => \N__36206\,
            I => \N__36154\
        );

    \I__6788\ : InMux
    port map (
            O => \N__36205\,
            I => \N__36145\
        );

    \I__6787\ : InMux
    port map (
            O => \N__36204\,
            I => \N__36145\
        );

    \I__6786\ : InMux
    port map (
            O => \N__36203\,
            I => \N__36145\
        );

    \I__6785\ : InMux
    port map (
            O => \N__36202\,
            I => \N__36145\
        );

    \I__6784\ : InMux
    port map (
            O => \N__36201\,
            I => \N__36134\
        );

    \I__6783\ : InMux
    port map (
            O => \N__36200\,
            I => \N__36134\
        );

    \I__6782\ : InMux
    port map (
            O => \N__36199\,
            I => \N__36134\
        );

    \I__6781\ : InMux
    port map (
            O => \N__36198\,
            I => \N__36134\
        );

    \I__6780\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36134\
        );

    \I__6779\ : InMux
    port map (
            O => \N__36196\,
            I => \N__36125\
        );

    \I__6778\ : InMux
    port map (
            O => \N__36195\,
            I => \N__36125\
        );

    \I__6777\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36125\
        );

    \I__6776\ : InMux
    port map (
            O => \N__36193\,
            I => \N__36125\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__36184\,
            I => \N__36114\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__36175\,
            I => \N__36114\
        );

    \I__6773\ : Span4Mux_v
    port map (
            O => \N__36172\,
            I => \N__36114\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__36163\,
            I => \N__36114\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__36154\,
            I => \N__36114\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__36145\,
            I => \N__36109\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__36134\,
            I => \N__36109\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__36125\,
            I => \phase_controller_inst2.stoper_hc.start_latched_i_0\
        );

    \I__6767\ : Odrv4
    port map (
            O => \N__36114\,
            I => \phase_controller_inst2.stoper_hc.start_latched_i_0\
        );

    \I__6766\ : Odrv12
    port map (
            O => \N__36109\,
            I => \phase_controller_inst2.stoper_hc.start_latched_i_0\
        );

    \I__6765\ : InMux
    port map (
            O => \N__36102\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_30\
        );

    \I__6764\ : InMux
    port map (
            O => \N__36099\,
            I => \N__36094\
        );

    \I__6763\ : InMux
    port map (
            O => \N__36098\,
            I => \N__36089\
        );

    \I__6762\ : InMux
    port map (
            O => \N__36097\,
            I => \N__36089\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__36094\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_31\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__36089\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_31\
        );

    \I__6759\ : CEMux
    port map (
            O => \N__36084\,
            I => \N__36081\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__36081\,
            I => \N__36078\
        );

    \I__6757\ : Span4Mux_v
    port map (
            O => \N__36078\,
            I => \N__36073\
        );

    \I__6756\ : CEMux
    port map (
            O => \N__36077\,
            I => \N__36070\
        );

    \I__6755\ : CEMux
    port map (
            O => \N__36076\,
            I => \N__36067\
        );

    \I__6754\ : Span4Mux_v
    port map (
            O => \N__36073\,
            I => \N__36062\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__36070\,
            I => \N__36062\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__36067\,
            I => \N__36059\
        );

    \I__6751\ : Span4Mux_v
    port map (
            O => \N__36062\,
            I => \N__36055\
        );

    \I__6750\ : Span12Mux_h
    port map (
            O => \N__36059\,
            I => \N__36052\
        );

    \I__6749\ : CEMux
    port map (
            O => \N__36058\,
            I => \N__36049\
        );

    \I__6748\ : Odrv4
    port map (
            O => \N__36055\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__6747\ : Odrv12
    port map (
            O => \N__36052\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__36049\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__6745\ : InMux
    port map (
            O => \N__36042\,
            I => \N__36036\
        );

    \I__6744\ : InMux
    port map (
            O => \N__36041\,
            I => \N__36036\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__36036\,
            I => \N__36033\
        );

    \I__6742\ : Odrv4
    port map (
            O => \N__36033\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_22\
        );

    \I__6741\ : InMux
    port map (
            O => \N__36030\,
            I => \N__36026\
        );

    \I__6740\ : InMux
    port map (
            O => \N__36029\,
            I => \N__36023\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__36026\,
            I => \N__36020\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__36023\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26\
        );

    \I__6737\ : Odrv4
    port map (
            O => \N__36020\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26\
        );

    \I__6736\ : InMux
    port map (
            O => \N__36015\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_16\
        );

    \I__6735\ : InMux
    port map (
            O => \N__36012\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_17\
        );

    \I__6734\ : InMux
    port map (
            O => \N__36009\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_18\
        );

    \I__6733\ : InMux
    port map (
            O => \N__36006\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_19\
        );

    \I__6732\ : InMux
    port map (
            O => \N__36003\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_20\
        );

    \I__6731\ : InMux
    port map (
            O => \N__36000\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_21\
        );

    \I__6730\ : InMux
    port map (
            O => \N__35997\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_22\
        );

    \I__6729\ : InMux
    port map (
            O => \N__35994\,
            I => \bfn_13_10_0_\
        );

    \I__6728\ : InMux
    port map (
            O => \N__35991\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_24\
        );

    \I__6727\ : InMux
    port map (
            O => \N__35988\,
            I => \bfn_13_8_0_\
        );

    \I__6726\ : InMux
    port map (
            O => \N__35985\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_8\
        );

    \I__6725\ : InMux
    port map (
            O => \N__35982\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_9\
        );

    \I__6724\ : InMux
    port map (
            O => \N__35979\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_10\
        );

    \I__6723\ : InMux
    port map (
            O => \N__35976\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_11\
        );

    \I__6722\ : InMux
    port map (
            O => \N__35973\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_12\
        );

    \I__6721\ : InMux
    port map (
            O => \N__35970\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_13\
        );

    \I__6720\ : InMux
    port map (
            O => \N__35967\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_14\
        );

    \I__6719\ : InMux
    port map (
            O => \N__35964\,
            I => \bfn_13_9_0_\
        );

    \I__6718\ : InMux
    port map (
            O => \N__35961\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_0\
        );

    \I__6717\ : InMux
    port map (
            O => \N__35958\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_1\
        );

    \I__6716\ : InMux
    port map (
            O => \N__35955\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_2\
        );

    \I__6715\ : InMux
    port map (
            O => \N__35952\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_3\
        );

    \I__6714\ : InMux
    port map (
            O => \N__35949\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_4\
        );

    \I__6713\ : InMux
    port map (
            O => \N__35946\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_5\
        );

    \I__6712\ : InMux
    port map (
            O => \N__35943\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_6\
        );

    \I__6711\ : InMux
    port map (
            O => \N__35940\,
            I => \N__35935\
        );

    \I__6710\ : InMux
    port map (
            O => \N__35939\,
            I => \N__35930\
        );

    \I__6709\ : InMux
    port map (
            O => \N__35938\,
            I => \N__35930\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__35935\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_23\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__35930\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_23\
        );

    \I__6706\ : InMux
    port map (
            O => \N__35925\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_22\
        );

    \I__6705\ : InMux
    port map (
            O => \N__35922\,
            I => \N__35917\
        );

    \I__6704\ : InMux
    port map (
            O => \N__35921\,
            I => \N__35914\
        );

    \I__6703\ : InMux
    port map (
            O => \N__35920\,
            I => \N__35911\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__35917\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_24\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__35914\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_24\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__35911\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_24\
        );

    \I__6699\ : InMux
    port map (
            O => \N__35904\,
            I => \bfn_12_30_0_\
        );

    \I__6698\ : CascadeMux
    port map (
            O => \N__35901\,
            I => \N__35897\
        );

    \I__6697\ : InMux
    port map (
            O => \N__35900\,
            I => \N__35893\
        );

    \I__6696\ : InMux
    port map (
            O => \N__35897\,
            I => \N__35890\
        );

    \I__6695\ : InMux
    port map (
            O => \N__35896\,
            I => \N__35887\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__35893\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_25\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__35890\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_25\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__35887\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_25\
        );

    \I__6691\ : InMux
    port map (
            O => \N__35880\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_24\
        );

    \I__6690\ : CascadeMux
    port map (
            O => \N__35877\,
            I => \N__35873\
        );

    \I__6689\ : CascadeMux
    port map (
            O => \N__35876\,
            I => \N__35870\
        );

    \I__6688\ : InMux
    port map (
            O => \N__35873\,
            I => \N__35867\
        );

    \I__6687\ : InMux
    port map (
            O => \N__35870\,
            I => \N__35864\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__35867\,
            I => \N__35858\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__35864\,
            I => \N__35858\
        );

    \I__6684\ : InMux
    port map (
            O => \N__35863\,
            I => \N__35855\
        );

    \I__6683\ : Span4Mux_v
    port map (
            O => \N__35858\,
            I => \N__35852\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__35855\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_26\
        );

    \I__6681\ : Odrv4
    port map (
            O => \N__35852\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_26\
        );

    \I__6680\ : InMux
    port map (
            O => \N__35847\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_25\
        );

    \I__6679\ : InMux
    port map (
            O => \N__35844\,
            I => \N__35841\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__35841\,
            I => \N__35836\
        );

    \I__6677\ : InMux
    port map (
            O => \N__35840\,
            I => \N__35833\
        );

    \I__6676\ : InMux
    port map (
            O => \N__35839\,
            I => \N__35830\
        );

    \I__6675\ : Span4Mux_v
    port map (
            O => \N__35836\,
            I => \N__35827\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__35833\,
            I => \N__35824\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__35830\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_27\
        );

    \I__6672\ : Odrv4
    port map (
            O => \N__35827\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_27\
        );

    \I__6671\ : Odrv12
    port map (
            O => \N__35824\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_27\
        );

    \I__6670\ : InMux
    port map (
            O => \N__35817\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_26\
        );

    \I__6669\ : InMux
    port map (
            O => \N__35814\,
            I => \N__35810\
        );

    \I__6668\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35807\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__35810\,
            I => \N__35801\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__35807\,
            I => \N__35801\
        );

    \I__6665\ : InMux
    port map (
            O => \N__35806\,
            I => \N__35798\
        );

    \I__6664\ : Span4Mux_h
    port map (
            O => \N__35801\,
            I => \N__35795\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__35798\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_28\
        );

    \I__6662\ : Odrv4
    port map (
            O => \N__35795\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_28\
        );

    \I__6661\ : InMux
    port map (
            O => \N__35790\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_27\
        );

    \I__6660\ : InMux
    port map (
            O => \N__35787\,
            I => \N__35783\
        );

    \I__6659\ : InMux
    port map (
            O => \N__35786\,
            I => \N__35779\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__35783\,
            I => \N__35776\
        );

    \I__6657\ : InMux
    port map (
            O => \N__35782\,
            I => \N__35773\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__35779\,
            I => \N__35770\
        );

    \I__6655\ : Span4Mux_h
    port map (
            O => \N__35776\,
            I => \N__35767\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__35773\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_29\
        );

    \I__6653\ : Odrv4
    port map (
            O => \N__35770\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_29\
        );

    \I__6652\ : Odrv4
    port map (
            O => \N__35767\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_29\
        );

    \I__6651\ : InMux
    port map (
            O => \N__35760\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_28\
        );

    \I__6650\ : InMux
    port map (
            O => \N__35757\,
            I => \N__35752\
        );

    \I__6649\ : InMux
    port map (
            O => \N__35756\,
            I => \N__35749\
        );

    \I__6648\ : InMux
    port map (
            O => \N__35755\,
            I => \N__35746\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__35752\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_30\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__35749\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_30\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__35746\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_30\
        );

    \I__6644\ : InMux
    port map (
            O => \N__35739\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_29\
        );

    \I__6643\ : InMux
    port map (
            O => \N__35736\,
            I => \N__35696\
        );

    \I__6642\ : InMux
    port map (
            O => \N__35735\,
            I => \N__35696\
        );

    \I__6641\ : InMux
    port map (
            O => \N__35734\,
            I => \N__35696\
        );

    \I__6640\ : InMux
    port map (
            O => \N__35733\,
            I => \N__35696\
        );

    \I__6639\ : InMux
    port map (
            O => \N__35732\,
            I => \N__35689\
        );

    \I__6638\ : InMux
    port map (
            O => \N__35731\,
            I => \N__35689\
        );

    \I__6637\ : InMux
    port map (
            O => \N__35730\,
            I => \N__35689\
        );

    \I__6636\ : InMux
    port map (
            O => \N__35729\,
            I => \N__35680\
        );

    \I__6635\ : InMux
    port map (
            O => \N__35728\,
            I => \N__35680\
        );

    \I__6634\ : InMux
    port map (
            O => \N__35727\,
            I => \N__35680\
        );

    \I__6633\ : InMux
    port map (
            O => \N__35726\,
            I => \N__35680\
        );

    \I__6632\ : InMux
    port map (
            O => \N__35725\,
            I => \N__35669\
        );

    \I__6631\ : InMux
    port map (
            O => \N__35724\,
            I => \N__35669\
        );

    \I__6630\ : InMux
    port map (
            O => \N__35723\,
            I => \N__35669\
        );

    \I__6629\ : InMux
    port map (
            O => \N__35722\,
            I => \N__35669\
        );

    \I__6628\ : InMux
    port map (
            O => \N__35721\,
            I => \N__35669\
        );

    \I__6627\ : InMux
    port map (
            O => \N__35720\,
            I => \N__35660\
        );

    \I__6626\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35660\
        );

    \I__6625\ : InMux
    port map (
            O => \N__35718\,
            I => \N__35660\
        );

    \I__6624\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35660\
        );

    \I__6623\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35651\
        );

    \I__6622\ : InMux
    port map (
            O => \N__35715\,
            I => \N__35651\
        );

    \I__6621\ : InMux
    port map (
            O => \N__35714\,
            I => \N__35651\
        );

    \I__6620\ : InMux
    port map (
            O => \N__35713\,
            I => \N__35651\
        );

    \I__6619\ : InMux
    port map (
            O => \N__35712\,
            I => \N__35642\
        );

    \I__6618\ : InMux
    port map (
            O => \N__35711\,
            I => \N__35642\
        );

    \I__6617\ : InMux
    port map (
            O => \N__35710\,
            I => \N__35642\
        );

    \I__6616\ : InMux
    port map (
            O => \N__35709\,
            I => \N__35642\
        );

    \I__6615\ : InMux
    port map (
            O => \N__35708\,
            I => \N__35633\
        );

    \I__6614\ : InMux
    port map (
            O => \N__35707\,
            I => \N__35633\
        );

    \I__6613\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35633\
        );

    \I__6612\ : InMux
    port map (
            O => \N__35705\,
            I => \N__35633\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__35696\,
            I => \N__35630\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__35689\,
            I => \N__35627\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__35680\,
            I => \N__35616\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__35669\,
            I => \N__35616\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__35660\,
            I => \N__35616\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__35651\,
            I => \N__35616\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__35642\,
            I => \N__35616\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__35633\,
            I => \N__35613\
        );

    \I__6603\ : Span4Mux_h
    port map (
            O => \N__35630\,
            I => \N__35606\
        );

    \I__6602\ : Span4Mux_s3_v
    port map (
            O => \N__35627\,
            I => \N__35606\
        );

    \I__6601\ : Span4Mux_s3_v
    port map (
            O => \N__35616\,
            I => \N__35606\
        );

    \I__6600\ : Odrv12
    port map (
            O => \N__35613\,
            I => \phase_controller_inst1.stoper_tr.start_latched_i_0\
        );

    \I__6599\ : Odrv4
    port map (
            O => \N__35606\,
            I => \phase_controller_inst1.stoper_tr.start_latched_i_0\
        );

    \I__6598\ : InMux
    port map (
            O => \N__35601\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_30\
        );

    \I__6597\ : InMux
    port map (
            O => \N__35598\,
            I => \N__35593\
        );

    \I__6596\ : InMux
    port map (
            O => \N__35597\,
            I => \N__35590\
        );

    \I__6595\ : InMux
    port map (
            O => \N__35596\,
            I => \N__35587\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__35593\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_31\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__35590\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_31\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__35587\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_31\
        );

    \I__6591\ : CEMux
    port map (
            O => \N__35580\,
            I => \N__35568\
        );

    \I__6590\ : CEMux
    port map (
            O => \N__35579\,
            I => \N__35568\
        );

    \I__6589\ : CEMux
    port map (
            O => \N__35578\,
            I => \N__35568\
        );

    \I__6588\ : CEMux
    port map (
            O => \N__35577\,
            I => \N__35568\
        );

    \I__6587\ : GlobalMux
    port map (
            O => \N__35568\,
            I => \N__35565\
        );

    \I__6586\ : gio2CtrlBuf
    port map (
            O => \N__35565\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0_g\
        );

    \I__6585\ : InMux
    port map (
            O => \N__35562\,
            I => \N__35558\
        );

    \I__6584\ : InMux
    port map (
            O => \N__35561\,
            I => \N__35555\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__35558\,
            I => \N__35552\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__35555\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_15\
        );

    \I__6581\ : Odrv4
    port map (
            O => \N__35552\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_15\
        );

    \I__6580\ : InMux
    port map (
            O => \N__35547\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_14\
        );

    \I__6579\ : InMux
    port map (
            O => \N__35544\,
            I => \bfn_12_29_0_\
        );

    \I__6578\ : InMux
    port map (
            O => \N__35541\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_16\
        );

    \I__6577\ : InMux
    port map (
            O => \N__35538\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_17\
        );

    \I__6576\ : InMux
    port map (
            O => \N__35535\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_18\
        );

    \I__6575\ : InMux
    port map (
            O => \N__35532\,
            I => \N__35527\
        );

    \I__6574\ : InMux
    port map (
            O => \N__35531\,
            I => \N__35524\
        );

    \I__6573\ : InMux
    port map (
            O => \N__35530\,
            I => \N__35521\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__35527\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_20\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__35524\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_20\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__35521\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_20\
        );

    \I__6569\ : InMux
    port map (
            O => \N__35514\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_19\
        );

    \I__6568\ : CascadeMux
    port map (
            O => \N__35511\,
            I => \N__35507\
        );

    \I__6567\ : InMux
    port map (
            O => \N__35510\,
            I => \N__35503\
        );

    \I__6566\ : InMux
    port map (
            O => \N__35507\,
            I => \N__35500\
        );

    \I__6565\ : InMux
    port map (
            O => \N__35506\,
            I => \N__35497\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__35503\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_21\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__35500\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_21\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__35497\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_21\
        );

    \I__6561\ : InMux
    port map (
            O => \N__35490\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_20\
        );

    \I__6560\ : InMux
    port map (
            O => \N__35487\,
            I => \N__35482\
        );

    \I__6559\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35477\
        );

    \I__6558\ : InMux
    port map (
            O => \N__35485\,
            I => \N__35477\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__35482\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_22\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__35477\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_22\
        );

    \I__6555\ : InMux
    port map (
            O => \N__35472\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_21\
        );

    \I__6554\ : InMux
    port map (
            O => \N__35469\,
            I => \N__35465\
        );

    \I__6553\ : InMux
    port map (
            O => \N__35468\,
            I => \N__35462\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__35465\,
            I => \N__35459\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__35462\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_6\
        );

    \I__6550\ : Odrv4
    port map (
            O => \N__35459\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_6\
        );

    \I__6549\ : InMux
    port map (
            O => \N__35454\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_5\
        );

    \I__6548\ : InMux
    port map (
            O => \N__35451\,
            I => \N__35447\
        );

    \I__6547\ : InMux
    port map (
            O => \N__35450\,
            I => \N__35444\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__35447\,
            I => \N__35441\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__35444\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_7\
        );

    \I__6544\ : Odrv4
    port map (
            O => \N__35441\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_7\
        );

    \I__6543\ : InMux
    port map (
            O => \N__35436\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_6\
        );

    \I__6542\ : InMux
    port map (
            O => \N__35433\,
            I => \N__35429\
        );

    \I__6541\ : InMux
    port map (
            O => \N__35432\,
            I => \N__35426\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__35429\,
            I => \N__35423\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__35426\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_8\
        );

    \I__6538\ : Odrv4
    port map (
            O => \N__35423\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_8\
        );

    \I__6537\ : InMux
    port map (
            O => \N__35418\,
            I => \bfn_12_28_0_\
        );

    \I__6536\ : InMux
    port map (
            O => \N__35415\,
            I => \N__35411\
        );

    \I__6535\ : InMux
    port map (
            O => \N__35414\,
            I => \N__35408\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__35411\,
            I => \N__35405\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__35408\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_9\
        );

    \I__6532\ : Odrv4
    port map (
            O => \N__35405\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_9\
        );

    \I__6531\ : InMux
    port map (
            O => \N__35400\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_8\
        );

    \I__6530\ : InMux
    port map (
            O => \N__35397\,
            I => \N__35393\
        );

    \I__6529\ : InMux
    port map (
            O => \N__35396\,
            I => \N__35390\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__35393\,
            I => \N__35387\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__35390\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_10\
        );

    \I__6526\ : Odrv4
    port map (
            O => \N__35387\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_10\
        );

    \I__6525\ : InMux
    port map (
            O => \N__35382\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_9\
        );

    \I__6524\ : InMux
    port map (
            O => \N__35379\,
            I => \N__35375\
        );

    \I__6523\ : InMux
    port map (
            O => \N__35378\,
            I => \N__35372\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__35375\,
            I => \N__35369\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__35372\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_11\
        );

    \I__6520\ : Odrv4
    port map (
            O => \N__35369\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_11\
        );

    \I__6519\ : InMux
    port map (
            O => \N__35364\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_10\
        );

    \I__6518\ : InMux
    port map (
            O => \N__35361\,
            I => \N__35357\
        );

    \I__6517\ : InMux
    port map (
            O => \N__35360\,
            I => \N__35354\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__35357\,
            I => \N__35351\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__35354\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_12\
        );

    \I__6514\ : Odrv4
    port map (
            O => \N__35351\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_12\
        );

    \I__6513\ : InMux
    port map (
            O => \N__35346\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_11\
        );

    \I__6512\ : InMux
    port map (
            O => \N__35343\,
            I => \N__35339\
        );

    \I__6511\ : InMux
    port map (
            O => \N__35342\,
            I => \N__35336\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__35339\,
            I => \N__35333\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__35336\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_13\
        );

    \I__6508\ : Odrv4
    port map (
            O => \N__35333\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_13\
        );

    \I__6507\ : InMux
    port map (
            O => \N__35328\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_12\
        );

    \I__6506\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35321\
        );

    \I__6505\ : InMux
    port map (
            O => \N__35324\,
            I => \N__35318\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__35321\,
            I => \N__35315\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__35318\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_14\
        );

    \I__6502\ : Odrv4
    port map (
            O => \N__35315\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_14\
        );

    \I__6501\ : InMux
    port map (
            O => \N__35310\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_13\
        );

    \I__6500\ : InMux
    port map (
            O => \N__35307\,
            I => \N__35304\
        );

    \I__6499\ : LocalMux
    port map (
            O => \N__35304\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_4\
        );

    \I__6498\ : InMux
    port map (
            O => \N__35301\,
            I => \N__35297\
        );

    \I__6497\ : InMux
    port map (
            O => \N__35300\,
            I => \N__35294\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__35297\,
            I => \N__35291\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__35294\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26\
        );

    \I__6494\ : Odrv4
    port map (
            O => \N__35291\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26\
        );

    \I__6493\ : InMux
    port map (
            O => \N__35286\,
            I => \N__35282\
        );

    \I__6492\ : InMux
    port map (
            O => \N__35285\,
            I => \N__35279\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__35282\,
            I => \N__35276\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__35279\,
            I => \N__35273\
        );

    \I__6489\ : Odrv4
    port map (
            O => \N__35276\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27\
        );

    \I__6488\ : Odrv12
    port map (
            O => \N__35273\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27\
        );

    \I__6487\ : InMux
    port map (
            O => \N__35268\,
            I => \N__35265\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__35265\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26\
        );

    \I__6485\ : CascadeMux
    port map (
            O => \N__35262\,
            I => \N__35258\
        );

    \I__6484\ : InMux
    port map (
            O => \N__35261\,
            I => \N__35255\
        );

    \I__6483\ : InMux
    port map (
            O => \N__35258\,
            I => \N__35252\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__35255\,
            I => \phase_controller_inst1.stoper_tr.counter\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__35252\,
            I => \phase_controller_inst1.stoper_tr.counter\
        );

    \I__6480\ : InMux
    port map (
            O => \N__35247\,
            I => \N__35243\
        );

    \I__6479\ : InMux
    port map (
            O => \N__35246\,
            I => \N__35240\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__35243\,
            I => \N__35237\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__35240\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_0\
        );

    \I__6476\ : Odrv4
    port map (
            O => \N__35237\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_0\
        );

    \I__6475\ : InMux
    port map (
            O => \N__35232\,
            I => \N__35228\
        );

    \I__6474\ : InMux
    port map (
            O => \N__35231\,
            I => \N__35225\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__35228\,
            I => \N__35222\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__35225\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_1\
        );

    \I__6471\ : Odrv4
    port map (
            O => \N__35222\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_1\
        );

    \I__6470\ : InMux
    port map (
            O => \N__35217\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_0\
        );

    \I__6469\ : InMux
    port map (
            O => \N__35214\,
            I => \N__35211\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__35211\,
            I => \N__35207\
        );

    \I__6467\ : InMux
    port map (
            O => \N__35210\,
            I => \N__35204\
        );

    \I__6466\ : Span12Mux_h
    port map (
            O => \N__35207\,
            I => \N__35201\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__35204\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_2\
        );

    \I__6464\ : Odrv12
    port map (
            O => \N__35201\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_2\
        );

    \I__6463\ : InMux
    port map (
            O => \N__35196\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_1\
        );

    \I__6462\ : InMux
    port map (
            O => \N__35193\,
            I => \N__35190\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__35190\,
            I => \N__35186\
        );

    \I__6460\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35183\
        );

    \I__6459\ : Span4Mux_v
    port map (
            O => \N__35186\,
            I => \N__35180\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__35183\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_3\
        );

    \I__6457\ : Odrv4
    port map (
            O => \N__35180\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_3\
        );

    \I__6456\ : InMux
    port map (
            O => \N__35175\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_2\
        );

    \I__6455\ : InMux
    port map (
            O => \N__35172\,
            I => \N__35168\
        );

    \I__6454\ : InMux
    port map (
            O => \N__35171\,
            I => \N__35165\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__35168\,
            I => \N__35162\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__35165\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_4\
        );

    \I__6451\ : Odrv4
    port map (
            O => \N__35162\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_4\
        );

    \I__6450\ : InMux
    port map (
            O => \N__35157\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_3\
        );

    \I__6449\ : InMux
    port map (
            O => \N__35154\,
            I => \N__35151\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__35151\,
            I => \N__35147\
        );

    \I__6447\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35144\
        );

    \I__6446\ : Span4Mux_h
    port map (
            O => \N__35147\,
            I => \N__35141\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__35144\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_5\
        );

    \I__6444\ : Odrv4
    port map (
            O => \N__35141\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_5\
        );

    \I__6443\ : InMux
    port map (
            O => \N__35136\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_4\
        );

    \I__6442\ : InMux
    port map (
            O => \N__35133\,
            I => \N__35129\
        );

    \I__6441\ : InMux
    port map (
            O => \N__35132\,
            I => \N__35126\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__35129\,
            I => \N__35121\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__35126\,
            I => \N__35121\
        );

    \I__6438\ : Span4Mux_v
    port map (
            O => \N__35121\,
            I => \N__35118\
        );

    \I__6437\ : Odrv4
    port map (
            O => \N__35118\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_24\
        );

    \I__6436\ : CascadeMux
    port map (
            O => \N__35115\,
            I => \N__35111\
        );

    \I__6435\ : InMux
    port map (
            O => \N__35114\,
            I => \N__35108\
        );

    \I__6434\ : InMux
    port map (
            O => \N__35111\,
            I => \N__35105\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__35108\,
            I => \N__35100\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__35105\,
            I => \N__35100\
        );

    \I__6431\ : Span4Mux_v
    port map (
            O => \N__35100\,
            I => \N__35097\
        );

    \I__6430\ : Odrv4
    port map (
            O => \N__35097\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20\
        );

    \I__6429\ : InMux
    port map (
            O => \N__35094\,
            I => \N__35091\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__35091\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_5\
        );

    \I__6427\ : InMux
    port map (
            O => \N__35088\,
            I => \N__35085\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__35085\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_3\
        );

    \I__6425\ : InMux
    port map (
            O => \N__35082\,
            I => \N__35079\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__35079\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ1Z_1\
        );

    \I__6423\ : InMux
    port map (
            O => \N__35076\,
            I => \N__35073\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__35073\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_2\
        );

    \I__6421\ : InMux
    port map (
            O => \N__35070\,
            I => \N__35067\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__35067\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_6\
        );

    \I__6419\ : InMux
    port map (
            O => \N__35064\,
            I => \N__35061\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__35061\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_8\
        );

    \I__6417\ : InMux
    port map (
            O => \N__35058\,
            I => \N__35055\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__35055\,
            I => \N__35052\
        );

    \I__6415\ : Span4Mux_v
    port map (
            O => \N__35052\,
            I => \N__35049\
        );

    \I__6414\ : Span4Mux_v
    port map (
            O => \N__35049\,
            I => \N__35046\
        );

    \I__6413\ : Odrv4
    port map (
            O => \N__35046\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_13\
        );

    \I__6412\ : CascadeMux
    port map (
            O => \N__35043\,
            I => \N__35039\
        );

    \I__6411\ : CascadeMux
    port map (
            O => \N__35042\,
            I => \N__35036\
        );

    \I__6410\ : InMux
    port map (
            O => \N__35039\,
            I => \N__35031\
        );

    \I__6409\ : InMux
    port map (
            O => \N__35036\,
            I => \N__35031\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__35031\,
            I => \N__35028\
        );

    \I__6407\ : Span4Mux_v
    port map (
            O => \N__35028\,
            I => \N__35025\
        );

    \I__6406\ : Span4Mux_h
    port map (
            O => \N__35025\,
            I => \N__35022\
        );

    \I__6405\ : Odrv4
    port map (
            O => \N__35022\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_23\
        );

    \I__6404\ : InMux
    port map (
            O => \N__35019\,
            I => \N__35016\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__35016\,
            I => \N__35013\
        );

    \I__6402\ : Span4Mux_v
    port map (
            O => \N__35013\,
            I => \N__35010\
        );

    \I__6401\ : Odrv4
    port map (
            O => \N__35010\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_9\
        );

    \I__6400\ : InMux
    port map (
            O => \N__35007\,
            I => \N__35003\
        );

    \I__6399\ : InMux
    port map (
            O => \N__35006\,
            I => \N__35000\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__35003\,
            I => \N__34997\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__35000\,
            I => \N__34994\
        );

    \I__6396\ : Span4Mux_v
    port map (
            O => \N__34997\,
            I => \N__34989\
        );

    \I__6395\ : Span4Mux_v
    port map (
            O => \N__34994\,
            I => \N__34989\
        );

    \I__6394\ : Odrv4
    port map (
            O => \N__34989\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21\
        );

    \I__6393\ : CascadeMux
    port map (
            O => \N__34986\,
            I => \N__34983\
        );

    \I__6392\ : InMux
    port map (
            O => \N__34983\,
            I => \N__34980\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__34980\,
            I => \N__34977\
        );

    \I__6390\ : Span4Mux_v
    port map (
            O => \N__34977\,
            I => \N__34974\
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__34974\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_0\
        );

    \I__6388\ : CascadeMux
    port map (
            O => \N__34971\,
            I => \N__34967\
        );

    \I__6387\ : InMux
    port map (
            O => \N__34970\,
            I => \N__34964\
        );

    \I__6386\ : InMux
    port map (
            O => \N__34967\,
            I => \N__34961\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__34964\,
            I => \N__34956\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__34961\,
            I => \N__34956\
        );

    \I__6383\ : Span4Mux_v
    port map (
            O => \N__34956\,
            I => \N__34953\
        );

    \I__6382\ : Odrv4
    port map (
            O => \N__34953\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25\
        );

    \I__6381\ : InMux
    port map (
            O => \N__34950\,
            I => \N__34946\
        );

    \I__6380\ : CascadeMux
    port map (
            O => \N__34949\,
            I => \N__34941\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__34946\,
            I => \N__34938\
        );

    \I__6378\ : InMux
    port map (
            O => \N__34945\,
            I => \N__34935\
        );

    \I__6377\ : InMux
    port map (
            O => \N__34944\,
            I => \N__34932\
        );

    \I__6376\ : InMux
    port map (
            O => \N__34941\,
            I => \N__34929\
        );

    \I__6375\ : Span4Mux_h
    port map (
            O => \N__34938\,
            I => \N__34926\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__34935\,
            I => \N__34919\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__34932\,
            I => \N__34919\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__34929\,
            I => \N__34919\
        );

    \I__6371\ : Span4Mux_v
    port map (
            O => \N__34926\,
            I => \N__34916\
        );

    \I__6370\ : Span4Mux_v
    port map (
            O => \N__34919\,
            I => \N__34913\
        );

    \I__6369\ : Odrv4
    port map (
            O => \N__34916\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28\
        );

    \I__6368\ : Odrv4
    port map (
            O => \N__34913\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28\
        );

    \I__6367\ : CascadeMux
    port map (
            O => \N__34908\,
            I => \N__34894\
        );

    \I__6366\ : InMux
    port map (
            O => \N__34907\,
            I => \N__34888\
        );

    \I__6365\ : InMux
    port map (
            O => \N__34906\,
            I => \N__34888\
        );

    \I__6364\ : CascadeMux
    port map (
            O => \N__34905\,
            I => \N__34884\
        );

    \I__6363\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34871\
        );

    \I__6362\ : InMux
    port map (
            O => \N__34903\,
            I => \N__34871\
        );

    \I__6361\ : InMux
    port map (
            O => \N__34902\,
            I => \N__34871\
        );

    \I__6360\ : InMux
    port map (
            O => \N__34901\,
            I => \N__34871\
        );

    \I__6359\ : InMux
    port map (
            O => \N__34900\,
            I => \N__34871\
        );

    \I__6358\ : InMux
    port map (
            O => \N__34899\,
            I => \N__34871\
        );

    \I__6357\ : InMux
    port map (
            O => \N__34898\,
            I => \N__34866\
        );

    \I__6356\ : InMux
    port map (
            O => \N__34897\,
            I => \N__34866\
        );

    \I__6355\ : InMux
    port map (
            O => \N__34894\,
            I => \N__34861\
        );

    \I__6354\ : InMux
    port map (
            O => \N__34893\,
            I => \N__34861\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__34888\,
            I => \N__34840\
        );

    \I__6352\ : InMux
    port map (
            O => \N__34887\,
            I => \N__34835\
        );

    \I__6351\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34835\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__34871\,
            I => \N__34832\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__34866\,
            I => \N__34827\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__34861\,
            I => \N__34827\
        );

    \I__6347\ : CascadeMux
    port map (
            O => \N__34860\,
            I => \N__34824\
        );

    \I__6346\ : CascadeMux
    port map (
            O => \N__34859\,
            I => \N__34821\
        );

    \I__6345\ : InMux
    port map (
            O => \N__34858\,
            I => \N__34818\
        );

    \I__6344\ : InMux
    port map (
            O => \N__34857\,
            I => \N__34811\
        );

    \I__6343\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34811\
        );

    \I__6342\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34811\
        );

    \I__6341\ : CascadeMux
    port map (
            O => \N__34854\,
            I => \N__34804\
        );

    \I__6340\ : CascadeMux
    port map (
            O => \N__34853\,
            I => \N__34801\
        );

    \I__6339\ : CascadeMux
    port map (
            O => \N__34852\,
            I => \N__34794\
        );

    \I__6338\ : CascadeMux
    port map (
            O => \N__34851\,
            I => \N__34788\
        );

    \I__6337\ : CascadeMux
    port map (
            O => \N__34850\,
            I => \N__34779\
        );

    \I__6336\ : CascadeMux
    port map (
            O => \N__34849\,
            I => \N__34776\
        );

    \I__6335\ : CascadeMux
    port map (
            O => \N__34848\,
            I => \N__34769\
        );

    \I__6334\ : CascadeMux
    port map (
            O => \N__34847\,
            I => \N__34766\
        );

    \I__6333\ : CascadeMux
    port map (
            O => \N__34846\,
            I => \N__34759\
        );

    \I__6332\ : CascadeMux
    port map (
            O => \N__34845\,
            I => \N__34755\
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__34844\,
            I => \N__34751\
        );

    \I__6330\ : CascadeMux
    port map (
            O => \N__34843\,
            I => \N__34747\
        );

    \I__6329\ : Span4Mux_h
    port map (
            O => \N__34840\,
            I => \N__34726\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__34835\,
            I => \N__34726\
        );

    \I__6327\ : Span4Mux_h
    port map (
            O => \N__34832\,
            I => \N__34726\
        );

    \I__6326\ : Span4Mux_v
    port map (
            O => \N__34827\,
            I => \N__34723\
        );

    \I__6325\ : InMux
    port map (
            O => \N__34824\,
            I => \N__34720\
        );

    \I__6324\ : InMux
    port map (
            O => \N__34821\,
            I => \N__34717\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__34818\,
            I => \N__34712\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__34811\,
            I => \N__34712\
        );

    \I__6321\ : InMux
    port map (
            O => \N__34810\,
            I => \N__34703\
        );

    \I__6320\ : InMux
    port map (
            O => \N__34809\,
            I => \N__34703\
        );

    \I__6319\ : InMux
    port map (
            O => \N__34808\,
            I => \N__34703\
        );

    \I__6318\ : InMux
    port map (
            O => \N__34807\,
            I => \N__34703\
        );

    \I__6317\ : InMux
    port map (
            O => \N__34804\,
            I => \N__34700\
        );

    \I__6316\ : InMux
    port map (
            O => \N__34801\,
            I => \N__34697\
        );

    \I__6315\ : InMux
    port map (
            O => \N__34800\,
            I => \N__34686\
        );

    \I__6314\ : InMux
    port map (
            O => \N__34799\,
            I => \N__34686\
        );

    \I__6313\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34686\
        );

    \I__6312\ : InMux
    port map (
            O => \N__34797\,
            I => \N__34686\
        );

    \I__6311\ : InMux
    port map (
            O => \N__34794\,
            I => \N__34686\
        );

    \I__6310\ : CascadeMux
    port map (
            O => \N__34793\,
            I => \N__34678\
        );

    \I__6309\ : CascadeMux
    port map (
            O => \N__34792\,
            I => \N__34673\
        );

    \I__6308\ : CascadeMux
    port map (
            O => \N__34791\,
            I => \N__34670\
        );

    \I__6307\ : InMux
    port map (
            O => \N__34788\,
            I => \N__34667\
        );

    \I__6306\ : InMux
    port map (
            O => \N__34787\,
            I => \N__34664\
        );

    \I__6305\ : CascadeMux
    port map (
            O => \N__34786\,
            I => \N__34661\
        );

    \I__6304\ : CascadeMux
    port map (
            O => \N__34785\,
            I => \N__34658\
        );

    \I__6303\ : InMux
    port map (
            O => \N__34784\,
            I => \N__34647\
        );

    \I__6302\ : InMux
    port map (
            O => \N__34783\,
            I => \N__34647\
        );

    \I__6301\ : InMux
    port map (
            O => \N__34782\,
            I => \N__34647\
        );

    \I__6300\ : InMux
    port map (
            O => \N__34779\,
            I => \N__34647\
        );

    \I__6299\ : InMux
    port map (
            O => \N__34776\,
            I => \N__34647\
        );

    \I__6298\ : InMux
    port map (
            O => \N__34775\,
            I => \N__34644\
        );

    \I__6297\ : InMux
    port map (
            O => \N__34774\,
            I => \N__34630\
        );

    \I__6296\ : InMux
    port map (
            O => \N__34773\,
            I => \N__34630\
        );

    \I__6295\ : InMux
    port map (
            O => \N__34772\,
            I => \N__34630\
        );

    \I__6294\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34625\
        );

    \I__6293\ : InMux
    port map (
            O => \N__34766\,
            I => \N__34625\
        );

    \I__6292\ : CascadeMux
    port map (
            O => \N__34765\,
            I => \N__34622\
        );

    \I__6291\ : CascadeMux
    port map (
            O => \N__34764\,
            I => \N__34618\
        );

    \I__6290\ : CascadeMux
    port map (
            O => \N__34763\,
            I => \N__34614\
        );

    \I__6289\ : InMux
    port map (
            O => \N__34762\,
            I => \N__34596\
        );

    \I__6288\ : InMux
    port map (
            O => \N__34759\,
            I => \N__34596\
        );

    \I__6287\ : InMux
    port map (
            O => \N__34758\,
            I => \N__34596\
        );

    \I__6286\ : InMux
    port map (
            O => \N__34755\,
            I => \N__34596\
        );

    \I__6285\ : InMux
    port map (
            O => \N__34754\,
            I => \N__34596\
        );

    \I__6284\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34596\
        );

    \I__6283\ : InMux
    port map (
            O => \N__34750\,
            I => \N__34596\
        );

    \I__6282\ : InMux
    port map (
            O => \N__34747\,
            I => \N__34596\
        );

    \I__6281\ : CascadeMux
    port map (
            O => \N__34746\,
            I => \N__34593\
        );

    \I__6280\ : CascadeMux
    port map (
            O => \N__34745\,
            I => \N__34589\
        );

    \I__6279\ : CascadeMux
    port map (
            O => \N__34744\,
            I => \N__34585\
        );

    \I__6278\ : CascadeMux
    port map (
            O => \N__34743\,
            I => \N__34581\
        );

    \I__6277\ : CascadeMux
    port map (
            O => \N__34742\,
            I => \N__34577\
        );

    \I__6276\ : CascadeMux
    port map (
            O => \N__34741\,
            I => \N__34573\
        );

    \I__6275\ : CascadeMux
    port map (
            O => \N__34740\,
            I => \N__34569\
        );

    \I__6274\ : CascadeMux
    port map (
            O => \N__34739\,
            I => \N__34565\
        );

    \I__6273\ : CascadeMux
    port map (
            O => \N__34738\,
            I => \N__34560\
        );

    \I__6272\ : CascadeMux
    port map (
            O => \N__34737\,
            I => \N__34556\
        );

    \I__6271\ : CascadeMux
    port map (
            O => \N__34736\,
            I => \N__34552\
        );

    \I__6270\ : CascadeMux
    port map (
            O => \N__34735\,
            I => \N__34547\
        );

    \I__6269\ : CascadeMux
    port map (
            O => \N__34734\,
            I => \N__34543\
        );

    \I__6268\ : CascadeMux
    port map (
            O => \N__34733\,
            I => \N__34539\
        );

    \I__6267\ : Span4Mux_v
    port map (
            O => \N__34726\,
            I => \N__34529\
        );

    \I__6266\ : Span4Mux_h
    port map (
            O => \N__34723\,
            I => \N__34529\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__34720\,
            I => \N__34529\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__34717\,
            I => \N__34529\
        );

    \I__6263\ : Span4Mux_v
    port map (
            O => \N__34712\,
            I => \N__34526\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__34703\,
            I => \N__34517\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__34700\,
            I => \N__34517\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__34697\,
            I => \N__34517\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__34686\,
            I => \N__34517\
        );

    \I__6258\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34508\
        );

    \I__6257\ : InMux
    port map (
            O => \N__34684\,
            I => \N__34508\
        );

    \I__6256\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34508\
        );

    \I__6255\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34508\
        );

    \I__6254\ : InMux
    port map (
            O => \N__34681\,
            I => \N__34505\
        );

    \I__6253\ : InMux
    port map (
            O => \N__34678\,
            I => \N__34494\
        );

    \I__6252\ : InMux
    port map (
            O => \N__34677\,
            I => \N__34494\
        );

    \I__6251\ : InMux
    port map (
            O => \N__34676\,
            I => \N__34494\
        );

    \I__6250\ : InMux
    port map (
            O => \N__34673\,
            I => \N__34494\
        );

    \I__6249\ : InMux
    port map (
            O => \N__34670\,
            I => \N__34494\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__34667\,
            I => \N__34485\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__34664\,
            I => \N__34485\
        );

    \I__6246\ : InMux
    port map (
            O => \N__34661\,
            I => \N__34482\
        );

    \I__6245\ : InMux
    port map (
            O => \N__34658\,
            I => \N__34479\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__34647\,
            I => \N__34474\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__34644\,
            I => \N__34474\
        );

    \I__6242\ : CascadeMux
    port map (
            O => \N__34643\,
            I => \N__34471\
        );

    \I__6241\ : CascadeMux
    port map (
            O => \N__34642\,
            I => \N__34467\
        );

    \I__6240\ : CascadeMux
    port map (
            O => \N__34641\,
            I => \N__34463\
        );

    \I__6239\ : CascadeMux
    port map (
            O => \N__34640\,
            I => \N__34459\
        );

    \I__6238\ : CascadeMux
    port map (
            O => \N__34639\,
            I => \N__34455\
        );

    \I__6237\ : CascadeMux
    port map (
            O => \N__34638\,
            I => \N__34451\
        );

    \I__6236\ : CascadeMux
    port map (
            O => \N__34637\,
            I => \N__34447\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__34630\,
            I => \N__34441\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__34625\,
            I => \N__34441\
        );

    \I__6233\ : InMux
    port map (
            O => \N__34622\,
            I => \N__34428\
        );

    \I__6232\ : InMux
    port map (
            O => \N__34621\,
            I => \N__34428\
        );

    \I__6231\ : InMux
    port map (
            O => \N__34618\,
            I => \N__34428\
        );

    \I__6230\ : InMux
    port map (
            O => \N__34617\,
            I => \N__34428\
        );

    \I__6229\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34428\
        );

    \I__6228\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34428\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__34596\,
            I => \N__34425\
        );

    \I__6226\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34408\
        );

    \I__6225\ : InMux
    port map (
            O => \N__34592\,
            I => \N__34408\
        );

    \I__6224\ : InMux
    port map (
            O => \N__34589\,
            I => \N__34408\
        );

    \I__6223\ : InMux
    port map (
            O => \N__34588\,
            I => \N__34408\
        );

    \I__6222\ : InMux
    port map (
            O => \N__34585\,
            I => \N__34408\
        );

    \I__6221\ : InMux
    port map (
            O => \N__34584\,
            I => \N__34408\
        );

    \I__6220\ : InMux
    port map (
            O => \N__34581\,
            I => \N__34408\
        );

    \I__6219\ : InMux
    port map (
            O => \N__34580\,
            I => \N__34408\
        );

    \I__6218\ : InMux
    port map (
            O => \N__34577\,
            I => \N__34391\
        );

    \I__6217\ : InMux
    port map (
            O => \N__34576\,
            I => \N__34391\
        );

    \I__6216\ : InMux
    port map (
            O => \N__34573\,
            I => \N__34391\
        );

    \I__6215\ : InMux
    port map (
            O => \N__34572\,
            I => \N__34391\
        );

    \I__6214\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34391\
        );

    \I__6213\ : InMux
    port map (
            O => \N__34568\,
            I => \N__34391\
        );

    \I__6212\ : InMux
    port map (
            O => \N__34565\,
            I => \N__34391\
        );

    \I__6211\ : InMux
    port map (
            O => \N__34564\,
            I => \N__34391\
        );

    \I__6210\ : InMux
    port map (
            O => \N__34563\,
            I => \N__34376\
        );

    \I__6209\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34376\
        );

    \I__6208\ : InMux
    port map (
            O => \N__34559\,
            I => \N__34376\
        );

    \I__6207\ : InMux
    port map (
            O => \N__34556\,
            I => \N__34376\
        );

    \I__6206\ : InMux
    port map (
            O => \N__34555\,
            I => \N__34376\
        );

    \I__6205\ : InMux
    port map (
            O => \N__34552\,
            I => \N__34376\
        );

    \I__6204\ : InMux
    port map (
            O => \N__34551\,
            I => \N__34376\
        );

    \I__6203\ : InMux
    port map (
            O => \N__34550\,
            I => \N__34373\
        );

    \I__6202\ : InMux
    port map (
            O => \N__34547\,
            I => \N__34360\
        );

    \I__6201\ : InMux
    port map (
            O => \N__34546\,
            I => \N__34360\
        );

    \I__6200\ : InMux
    port map (
            O => \N__34543\,
            I => \N__34360\
        );

    \I__6199\ : InMux
    port map (
            O => \N__34542\,
            I => \N__34360\
        );

    \I__6198\ : InMux
    port map (
            O => \N__34539\,
            I => \N__34360\
        );

    \I__6197\ : InMux
    port map (
            O => \N__34538\,
            I => \N__34360\
        );

    \I__6196\ : Span4Mux_v
    port map (
            O => \N__34529\,
            I => \N__34357\
        );

    \I__6195\ : Span4Mux_h
    port map (
            O => \N__34526\,
            I => \N__34346\
        );

    \I__6194\ : Span4Mux_v
    port map (
            O => \N__34517\,
            I => \N__34346\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__34508\,
            I => \N__34346\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34346\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__34494\,
            I => \N__34346\
        );

    \I__6190\ : InMux
    port map (
            O => \N__34493\,
            I => \N__34337\
        );

    \I__6189\ : InMux
    port map (
            O => \N__34492\,
            I => \N__34337\
        );

    \I__6188\ : InMux
    port map (
            O => \N__34491\,
            I => \N__34337\
        );

    \I__6187\ : InMux
    port map (
            O => \N__34490\,
            I => \N__34337\
        );

    \I__6186\ : Span4Mux_v
    port map (
            O => \N__34485\,
            I => \N__34328\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__34482\,
            I => \N__34328\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__34479\,
            I => \N__34328\
        );

    \I__6183\ : Span4Mux_h
    port map (
            O => \N__34474\,
            I => \N__34328\
        );

    \I__6182\ : InMux
    port map (
            O => \N__34471\,
            I => \N__34311\
        );

    \I__6181\ : InMux
    port map (
            O => \N__34470\,
            I => \N__34311\
        );

    \I__6180\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34311\
        );

    \I__6179\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34311\
        );

    \I__6178\ : InMux
    port map (
            O => \N__34463\,
            I => \N__34311\
        );

    \I__6177\ : InMux
    port map (
            O => \N__34462\,
            I => \N__34311\
        );

    \I__6176\ : InMux
    port map (
            O => \N__34459\,
            I => \N__34311\
        );

    \I__6175\ : InMux
    port map (
            O => \N__34458\,
            I => \N__34311\
        );

    \I__6174\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34298\
        );

    \I__6173\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34298\
        );

    \I__6172\ : InMux
    port map (
            O => \N__34451\,
            I => \N__34298\
        );

    \I__6171\ : InMux
    port map (
            O => \N__34450\,
            I => \N__34298\
        );

    \I__6170\ : InMux
    port map (
            O => \N__34447\,
            I => \N__34298\
        );

    \I__6169\ : InMux
    port map (
            O => \N__34446\,
            I => \N__34298\
        );

    \I__6168\ : Sp12to4
    port map (
            O => \N__34441\,
            I => \N__34281\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__34428\,
            I => \N__34281\
        );

    \I__6166\ : Span12Mux_s9_v
    port map (
            O => \N__34425\,
            I => \N__34281\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__34408\,
            I => \N__34281\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__34391\,
            I => \N__34281\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__34376\,
            I => \N__34281\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__34373\,
            I => \N__34281\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__34360\,
            I => \N__34281\
        );

    \I__6160\ : Odrv4
    port map (
            O => \N__34357\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6159\ : Odrv4
    port map (
            O => \N__34346\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__34337\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6157\ : Odrv4
    port map (
            O => \N__34328\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__34311\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__34298\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6154\ : Odrv12
    port map (
            O => \N__34281\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6153\ : CascadeMux
    port map (
            O => \N__34266\,
            I => \N__34261\
        );

    \I__6152\ : InMux
    port map (
            O => \N__34265\,
            I => \N__34255\
        );

    \I__6151\ : InMux
    port map (
            O => \N__34264\,
            I => \N__34247\
        );

    \I__6150\ : InMux
    port map (
            O => \N__34261\,
            I => \N__34247\
        );

    \I__6149\ : InMux
    port map (
            O => \N__34260\,
            I => \N__34247\
        );

    \I__6148\ : InMux
    port map (
            O => \N__34259\,
            I => \N__34239\
        );

    \I__6147\ : InMux
    port map (
            O => \N__34258\,
            I => \N__34231\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__34255\,
            I => \N__34226\
        );

    \I__6145\ : InMux
    port map (
            O => \N__34254\,
            I => \N__34223\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__34247\,
            I => \N__34220\
        );

    \I__6143\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34215\
        );

    \I__6142\ : InMux
    port map (
            O => \N__34245\,
            I => \N__34215\
        );

    \I__6141\ : InMux
    port map (
            O => \N__34244\,
            I => \N__34212\
        );

    \I__6140\ : InMux
    port map (
            O => \N__34243\,
            I => \N__34203\
        );

    \I__6139\ : InMux
    port map (
            O => \N__34242\,
            I => \N__34203\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__34239\,
            I => \N__34182\
        );

    \I__6137\ : InMux
    port map (
            O => \N__34238\,
            I => \N__34177\
        );

    \I__6136\ : InMux
    port map (
            O => \N__34237\,
            I => \N__34177\
        );

    \I__6135\ : InMux
    port map (
            O => \N__34236\,
            I => \N__34174\
        );

    \I__6134\ : InMux
    port map (
            O => \N__34235\,
            I => \N__34169\
        );

    \I__6133\ : InMux
    port map (
            O => \N__34234\,
            I => \N__34169\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__34231\,
            I => \N__34166\
        );

    \I__6131\ : InMux
    port map (
            O => \N__34230\,
            I => \N__34163\
        );

    \I__6130\ : InMux
    port map (
            O => \N__34229\,
            I => \N__34160\
        );

    \I__6129\ : Span4Mux_v
    port map (
            O => \N__34226\,
            I => \N__34153\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__34223\,
            I => \N__34153\
        );

    \I__6127\ : Span4Mux_h
    port map (
            O => \N__34220\,
            I => \N__34153\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__34215\,
            I => \N__34148\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__34212\,
            I => \N__34148\
        );

    \I__6124\ : InMux
    port map (
            O => \N__34211\,
            I => \N__34141\
        );

    \I__6123\ : InMux
    port map (
            O => \N__34210\,
            I => \N__34141\
        );

    \I__6122\ : InMux
    port map (
            O => \N__34209\,
            I => \N__34141\
        );

    \I__6121\ : InMux
    port map (
            O => \N__34208\,
            I => \N__34138\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__34203\,
            I => \N__34130\
        );

    \I__6119\ : InMux
    port map (
            O => \N__34202\,
            I => \N__34117\
        );

    \I__6118\ : InMux
    port map (
            O => \N__34201\,
            I => \N__34117\
        );

    \I__6117\ : InMux
    port map (
            O => \N__34200\,
            I => \N__34117\
        );

    \I__6116\ : InMux
    port map (
            O => \N__34199\,
            I => \N__34117\
        );

    \I__6115\ : InMux
    port map (
            O => \N__34198\,
            I => \N__34117\
        );

    \I__6114\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34117\
        );

    \I__6113\ : InMux
    port map (
            O => \N__34196\,
            I => \N__34100\
        );

    \I__6112\ : InMux
    port map (
            O => \N__34195\,
            I => \N__34100\
        );

    \I__6111\ : InMux
    port map (
            O => \N__34194\,
            I => \N__34100\
        );

    \I__6110\ : InMux
    port map (
            O => \N__34193\,
            I => \N__34100\
        );

    \I__6109\ : InMux
    port map (
            O => \N__34192\,
            I => \N__34100\
        );

    \I__6108\ : InMux
    port map (
            O => \N__34191\,
            I => \N__34100\
        );

    \I__6107\ : InMux
    port map (
            O => \N__34190\,
            I => \N__34100\
        );

    \I__6106\ : InMux
    port map (
            O => \N__34189\,
            I => \N__34100\
        );

    \I__6105\ : InMux
    port map (
            O => \N__34188\,
            I => \N__34091\
        );

    \I__6104\ : InMux
    port map (
            O => \N__34187\,
            I => \N__34091\
        );

    \I__6103\ : InMux
    port map (
            O => \N__34186\,
            I => \N__34091\
        );

    \I__6102\ : InMux
    port map (
            O => \N__34185\,
            I => \N__34091\
        );

    \I__6101\ : Span4Mux_v
    port map (
            O => \N__34182\,
            I => \N__34083\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__34177\,
            I => \N__34080\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__34174\,
            I => \N__34057\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__34169\,
            I => \N__34046\
        );

    \I__6097\ : Span4Mux_h
    port map (
            O => \N__34166\,
            I => \N__34046\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__34163\,
            I => \N__34046\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__34160\,
            I => \N__34046\
        );

    \I__6094\ : Span4Mux_v
    port map (
            O => \N__34153\,
            I => \N__34046\
        );

    \I__6093\ : Span4Mux_v
    port map (
            O => \N__34148\,
            I => \N__34039\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__34141\,
            I => \N__34039\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__34138\,
            I => \N__34039\
        );

    \I__6090\ : InMux
    port map (
            O => \N__34137\,
            I => \N__34034\
        );

    \I__6089\ : InMux
    port map (
            O => \N__34136\,
            I => \N__34034\
        );

    \I__6088\ : InMux
    port map (
            O => \N__34135\,
            I => \N__34027\
        );

    \I__6087\ : InMux
    port map (
            O => \N__34134\,
            I => \N__34027\
        );

    \I__6086\ : InMux
    port map (
            O => \N__34133\,
            I => \N__34027\
        );

    \I__6085\ : Span4Mux_h
    port map (
            O => \N__34130\,
            I => \N__34018\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__34117\,
            I => \N__34018\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__34100\,
            I => \N__34018\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__34091\,
            I => \N__34018\
        );

    \I__6081\ : InMux
    port map (
            O => \N__34090\,
            I => \N__34015\
        );

    \I__6080\ : InMux
    port map (
            O => \N__34089\,
            I => \N__34006\
        );

    \I__6079\ : InMux
    port map (
            O => \N__34088\,
            I => \N__34006\
        );

    \I__6078\ : InMux
    port map (
            O => \N__34087\,
            I => \N__34006\
        );

    \I__6077\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34006\
        );

    \I__6076\ : Span4Mux_h
    port map (
            O => \N__34083\,
            I => \N__34001\
        );

    \I__6075\ : Span4Mux_v
    port map (
            O => \N__34080\,
            I => \N__34001\
        );

    \I__6074\ : InMux
    port map (
            O => \N__34079\,
            I => \N__33998\
        );

    \I__6073\ : InMux
    port map (
            O => \N__34078\,
            I => \N__33985\
        );

    \I__6072\ : InMux
    port map (
            O => \N__34077\,
            I => \N__33985\
        );

    \I__6071\ : InMux
    port map (
            O => \N__34076\,
            I => \N__33985\
        );

    \I__6070\ : InMux
    port map (
            O => \N__34075\,
            I => \N__33985\
        );

    \I__6069\ : InMux
    port map (
            O => \N__34074\,
            I => \N__33985\
        );

    \I__6068\ : InMux
    port map (
            O => \N__34073\,
            I => \N__33985\
        );

    \I__6067\ : InMux
    port map (
            O => \N__34072\,
            I => \N__33974\
        );

    \I__6066\ : InMux
    port map (
            O => \N__34071\,
            I => \N__33974\
        );

    \I__6065\ : InMux
    port map (
            O => \N__34070\,
            I => \N__33974\
        );

    \I__6064\ : InMux
    port map (
            O => \N__34069\,
            I => \N__33974\
        );

    \I__6063\ : InMux
    port map (
            O => \N__34068\,
            I => \N__33974\
        );

    \I__6062\ : InMux
    port map (
            O => \N__34067\,
            I => \N__33961\
        );

    \I__6061\ : InMux
    port map (
            O => \N__34066\,
            I => \N__33961\
        );

    \I__6060\ : InMux
    port map (
            O => \N__34065\,
            I => \N__33961\
        );

    \I__6059\ : InMux
    port map (
            O => \N__34064\,
            I => \N__33961\
        );

    \I__6058\ : InMux
    port map (
            O => \N__34063\,
            I => \N__33961\
        );

    \I__6057\ : InMux
    port map (
            O => \N__34062\,
            I => \N__33961\
        );

    \I__6056\ : InMux
    port map (
            O => \N__34061\,
            I => \N__33956\
        );

    \I__6055\ : InMux
    port map (
            O => \N__34060\,
            I => \N__33956\
        );

    \I__6054\ : Span4Mux_h
    port map (
            O => \N__34057\,
            I => \N__33949\
        );

    \I__6053\ : Span4Mux_v
    port map (
            O => \N__34046\,
            I => \N__33949\
        );

    \I__6052\ : Span4Mux_v
    port map (
            O => \N__34039\,
            I => \N__33949\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__34034\,
            I => \N__33942\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__34027\,
            I => \N__33942\
        );

    \I__6049\ : Span4Mux_v
    port map (
            O => \N__34018\,
            I => \N__33942\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__34015\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__34006\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6046\ : Odrv4
    port map (
            O => \N__34001\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__33998\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__33985\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__33974\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__33961\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__33956\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__33949\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6039\ : Odrv4
    port map (
            O => \N__33942\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6038\ : CascadeMux
    port map (
            O => \N__33921\,
            I => \N__33918\
        );

    \I__6037\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33912\
        );

    \I__6036\ : InMux
    port map (
            O => \N__33917\,
            I => \N__33907\
        );

    \I__6035\ : InMux
    port map (
            O => \N__33916\,
            I => \N__33907\
        );

    \I__6034\ : InMux
    port map (
            O => \N__33915\,
            I => \N__33904\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__33912\,
            I => \N__33901\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__33907\,
            I => \N__33898\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__33904\,
            I => \N__33895\
        );

    \I__6030\ : Span4Mux_v
    port map (
            O => \N__33901\,
            I => \N__33892\
        );

    \I__6029\ : Span4Mux_v
    port map (
            O => \N__33898\,
            I => \N__33887\
        );

    \I__6028\ : Span4Mux_h
    port map (
            O => \N__33895\,
            I => \N__33887\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__33892\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__6026\ : Odrv4
    port map (
            O => \N__33887\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__6025\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33877\
        );

    \I__6024\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33872\
        );

    \I__6023\ : InMux
    port map (
            O => \N__33880\,
            I => \N__33872\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__33877\,
            I => \N__33869\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__33872\,
            I => \N__33866\
        );

    \I__6020\ : Odrv4
    port map (
            O => \N__33869\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__6019\ : Odrv4
    port map (
            O => \N__33866\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__6018\ : InMux
    port map (
            O => \N__33861\,
            I => \N__33858\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__33858\,
            I => \N__33855\
        );

    \I__6016\ : Span4Mux_h
    port map (
            O => \N__33855\,
            I => \N__33852\
        );

    \I__6015\ : Odrv4
    port map (
            O => \N__33852\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__6014\ : InMux
    port map (
            O => \N__33849\,
            I => \N__33846\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__33846\,
            I => \N__33843\
        );

    \I__6012\ : Sp12to4
    port map (
            O => \N__33843\,
            I => \N__33840\
        );

    \I__6011\ : Odrv12
    port map (
            O => \N__33840\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_15\
        );

    \I__6010\ : InMux
    port map (
            O => \N__33837\,
            I => \N__33834\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__33834\,
            I => \N__33831\
        );

    \I__6008\ : Span4Mux_v
    port map (
            O => \N__33831\,
            I => \N__33828\
        );

    \I__6007\ : Odrv4
    port map (
            O => \N__33828\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_10\
        );

    \I__6006\ : InMux
    port map (
            O => \N__33825\,
            I => \N__33822\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__33822\,
            I => \N__33819\
        );

    \I__6004\ : Span4Mux_v
    port map (
            O => \N__33819\,
            I => \N__33816\
        );

    \I__6003\ : Odrv4
    port map (
            O => \N__33816\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_12\
        );

    \I__6002\ : InMux
    port map (
            O => \N__33813\,
            I => \N__33810\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__33810\,
            I => \N__33807\
        );

    \I__6000\ : Span4Mux_v
    port map (
            O => \N__33807\,
            I => \N__33804\
        );

    \I__5999\ : Odrv4
    port map (
            O => \N__33804\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_7\
        );

    \I__5998\ : InMux
    port map (
            O => \N__33801\,
            I => \N__33798\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__33798\,
            I => \N__33795\
        );

    \I__5996\ : Span4Mux_v
    port map (
            O => \N__33795\,
            I => \N__33792\
        );

    \I__5995\ : Odrv4
    port map (
            O => \N__33792\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_11\
        );

    \I__5994\ : InMux
    port map (
            O => \N__33789\,
            I => \N__33786\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__33786\,
            I => \N__33783\
        );

    \I__5992\ : Span4Mux_v
    port map (
            O => \N__33783\,
            I => \N__33780\
        );

    \I__5991\ : Odrv4
    port map (
            O => \N__33780\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_14\
        );

    \I__5990\ : InMux
    port map (
            O => \N__33777\,
            I => \N__33771\
        );

    \I__5989\ : InMux
    port map (
            O => \N__33776\,
            I => \N__33771\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__33771\,
            I => \N__33768\
        );

    \I__5987\ : Span4Mux_h
    port map (
            O => \N__33768\,
            I => \N__33765\
        );

    \I__5986\ : Span4Mux_v
    port map (
            O => \N__33765\,
            I => \N__33762\
        );

    \I__5985\ : Odrv4
    port map (
            O => \N__33762\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_22\
        );

    \I__5984\ : CEMux
    port map (
            O => \N__33759\,
            I => \N__33735\
        );

    \I__5983\ : CEMux
    port map (
            O => \N__33758\,
            I => \N__33735\
        );

    \I__5982\ : CEMux
    port map (
            O => \N__33757\,
            I => \N__33735\
        );

    \I__5981\ : CEMux
    port map (
            O => \N__33756\,
            I => \N__33735\
        );

    \I__5980\ : CEMux
    port map (
            O => \N__33755\,
            I => \N__33735\
        );

    \I__5979\ : CEMux
    port map (
            O => \N__33754\,
            I => \N__33735\
        );

    \I__5978\ : CEMux
    port map (
            O => \N__33753\,
            I => \N__33735\
        );

    \I__5977\ : CEMux
    port map (
            O => \N__33752\,
            I => \N__33735\
        );

    \I__5976\ : GlobalMux
    port map (
            O => \N__33735\,
            I => \N__33732\
        );

    \I__5975\ : gio2CtrlBuf
    port map (
            O => \N__33732\,
            I => \current_shift_inst.timer_s1.N_153_i_g\
        );

    \I__5974\ : InMux
    port map (
            O => \N__33729\,
            I => \N__33726\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__33726\,
            I => \N__33723\
        );

    \I__5972\ : Span4Mux_v
    port map (
            O => \N__33723\,
            I => \N__33719\
        );

    \I__5971\ : InMux
    port map (
            O => \N__33722\,
            I => \N__33716\
        );

    \I__5970\ : Odrv4
    port map (
            O => \N__33719\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__33716\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__5968\ : CascadeMux
    port map (
            O => \N__33711\,
            I => \N__33708\
        );

    \I__5967\ : InMux
    port map (
            O => \N__33708\,
            I => \N__33705\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__33705\,
            I => \N__33702\
        );

    \I__5965\ : Span4Mux_v
    port map (
            O => \N__33702\,
            I => \N__33699\
        );

    \I__5964\ : Odrv4
    port map (
            O => \N__33699\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__5963\ : InMux
    port map (
            O => \N__33696\,
            I => \N__33693\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__33693\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__5961\ : CascadeMux
    port map (
            O => \N__33690\,
            I => \N__33686\
        );

    \I__5960\ : CascadeMux
    port map (
            O => \N__33689\,
            I => \N__33683\
        );

    \I__5959\ : InMux
    port map (
            O => \N__33686\,
            I => \N__33679\
        );

    \I__5958\ : InMux
    port map (
            O => \N__33683\,
            I => \N__33676\
        );

    \I__5957\ : InMux
    port map (
            O => \N__33682\,
            I => \N__33673\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__33679\,
            I => \N__33670\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__33676\,
            I => \N__33666\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__33673\,
            I => \N__33663\
        );

    \I__5953\ : Span4Mux_v
    port map (
            O => \N__33670\,
            I => \N__33660\
        );

    \I__5952\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33657\
        );

    \I__5951\ : Span4Mux_h
    port map (
            O => \N__33666\,
            I => \N__33652\
        );

    \I__5950\ : Span4Mux_v
    port map (
            O => \N__33663\,
            I => \N__33652\
        );

    \I__5949\ : Sp12to4
    port map (
            O => \N__33660\,
            I => \N__33647\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__33657\,
            I => \N__33647\
        );

    \I__5947\ : Odrv4
    port map (
            O => \N__33652\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__5946\ : Odrv12
    port map (
            O => \N__33647\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__5945\ : InMux
    port map (
            O => \N__33642\,
            I => \N__33639\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__33639\,
            I => \N__33634\
        );

    \I__5943\ : InMux
    port map (
            O => \N__33638\,
            I => \N__33631\
        );

    \I__5942\ : InMux
    port map (
            O => \N__33637\,
            I => \N__33628\
        );

    \I__5941\ : Span4Mux_h
    port map (
            O => \N__33634\,
            I => \N__33625\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__33631\,
            I => \N__33622\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__33628\,
            I => \N__33619\
        );

    \I__5938\ : Odrv4
    port map (
            O => \N__33625\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__5937\ : Odrv4
    port map (
            O => \N__33622\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__33619\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__5935\ : InMux
    port map (
            O => \N__33612\,
            I => \N__33609\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__33609\,
            I => \N__33606\
        );

    \I__5933\ : Span4Mux_h
    port map (
            O => \N__33606\,
            I => \N__33603\
        );

    \I__5932\ : Odrv4
    port map (
            O => \N__33603\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\
        );

    \I__5931\ : CascadeMux
    port map (
            O => \N__33600\,
            I => \N__33597\
        );

    \I__5930\ : InMux
    port map (
            O => \N__33597\,
            I => \N__33593\
        );

    \I__5929\ : CascadeMux
    port map (
            O => \N__33596\,
            I => \N__33590\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__33593\,
            I => \N__33585\
        );

    \I__5927\ : InMux
    port map (
            O => \N__33590\,
            I => \N__33582\
        );

    \I__5926\ : InMux
    port map (
            O => \N__33589\,
            I => \N__33579\
        );

    \I__5925\ : InMux
    port map (
            O => \N__33588\,
            I => \N__33576\
        );

    \I__5924\ : Span4Mux_v
    port map (
            O => \N__33585\,
            I => \N__33569\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__33582\,
            I => \N__33569\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__33579\,
            I => \N__33569\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__33576\,
            I => \N__33566\
        );

    \I__5920\ : Sp12to4
    port map (
            O => \N__33569\,
            I => \N__33563\
        );

    \I__5919\ : Span4Mux_h
    port map (
            O => \N__33566\,
            I => \N__33560\
        );

    \I__5918\ : Odrv12
    port map (
            O => \N__33563\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__5917\ : Odrv4
    port map (
            O => \N__33560\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__5916\ : InMux
    port map (
            O => \N__33555\,
            I => \N__33552\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__33552\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__5914\ : CascadeMux
    port map (
            O => \N__33549\,
            I => \N__33546\
        );

    \I__5913\ : InMux
    port map (
            O => \N__33546\,
            I => \N__33541\
        );

    \I__5912\ : InMux
    port map (
            O => \N__33545\,
            I => \N__33536\
        );

    \I__5911\ : InMux
    port map (
            O => \N__33544\,
            I => \N__33536\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__33541\,
            I => \N__33533\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__33536\,
            I => \N__33530\
        );

    \I__5908\ : Span4Mux_h
    port map (
            O => \N__33533\,
            I => \N__33526\
        );

    \I__5907\ : Span4Mux_v
    port map (
            O => \N__33530\,
            I => \N__33523\
        );

    \I__5906\ : InMux
    port map (
            O => \N__33529\,
            I => \N__33520\
        );

    \I__5905\ : Odrv4
    port map (
            O => \N__33526\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__5904\ : Odrv4
    port map (
            O => \N__33523\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__33520\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__5902\ : CascadeMux
    port map (
            O => \N__33513\,
            I => \N__33510\
        );

    \I__5901\ : InMux
    port map (
            O => \N__33510\,
            I => \N__33505\
        );

    \I__5900\ : InMux
    port map (
            O => \N__33509\,
            I => \N__33502\
        );

    \I__5899\ : InMux
    port map (
            O => \N__33508\,
            I => \N__33499\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__33505\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__33502\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__33499\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__5895\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33489\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__33489\,
            I => \N__33486\
        );

    \I__5893\ : Span4Mux_h
    port map (
            O => \N__33486\,
            I => \N__33483\
        );

    \I__5892\ : Odrv4
    port map (
            O => \N__33483\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__5891\ : InMux
    port map (
            O => \N__33480\,
            I => \N__33477\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__33477\,
            I => \N__33474\
        );

    \I__5889\ : Span4Mux_v
    port map (
            O => \N__33474\,
            I => \N__33471\
        );

    \I__5888\ : Odrv4
    port map (
            O => \N__33471\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_14\
        );

    \I__5887\ : ClkMux
    port map (
            O => \N__33468\,
            I => \N__33465\
        );

    \I__5886\ : GlobalMux
    port map (
            O => \N__33465\,
            I => \N__33462\
        );

    \I__5885\ : gio2CtrlBuf
    port map (
            O => \N__33462\,
            I => delay_tr_input_c_g
        );

    \I__5884\ : InMux
    port map (
            O => \N__33459\,
            I => \N__33456\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__33456\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__5882\ : CascadeMux
    port map (
            O => \N__33453\,
            I => \N__33449\
        );

    \I__5881\ : CascadeMux
    port map (
            O => \N__33452\,
            I => \N__33446\
        );

    \I__5880\ : InMux
    port map (
            O => \N__33449\,
            I => \N__33443\
        );

    \I__5879\ : InMux
    port map (
            O => \N__33446\,
            I => \N__33440\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__33443\,
            I => \N__33435\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__33440\,
            I => \N__33432\
        );

    \I__5876\ : InMux
    port map (
            O => \N__33439\,
            I => \N__33429\
        );

    \I__5875\ : InMux
    port map (
            O => \N__33438\,
            I => \N__33426\
        );

    \I__5874\ : Span12Mux_v
    port map (
            O => \N__33435\,
            I => \N__33423\
        );

    \I__5873\ : Span12Mux_h
    port map (
            O => \N__33432\,
            I => \N__33416\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__33429\,
            I => \N__33416\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__33426\,
            I => \N__33416\
        );

    \I__5870\ : Odrv12
    port map (
            O => \N__33423\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__5869\ : Odrv12
    port map (
            O => \N__33416\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__5868\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33406\
        );

    \I__5867\ : InMux
    port map (
            O => \N__33410\,
            I => \N__33403\
        );

    \I__5866\ : InMux
    port map (
            O => \N__33409\,
            I => \N__33400\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__33406\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__33403\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__33400\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__5862\ : CascadeMux
    port map (
            O => \N__33393\,
            I => \N__33390\
        );

    \I__5861\ : InMux
    port map (
            O => \N__33390\,
            I => \N__33387\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__33387\,
            I => \N__33384\
        );

    \I__5859\ : Span4Mux_v
    port map (
            O => \N__33384\,
            I => \N__33381\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__33381\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\
        );

    \I__5857\ : InMux
    port map (
            O => \N__33378\,
            I => \N__33375\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__33375\,
            I => \N__33371\
        );

    \I__5855\ : InMux
    port map (
            O => \N__33374\,
            I => \N__33368\
        );

    \I__5854\ : Span4Mux_h
    port map (
            O => \N__33371\,
            I => \N__33364\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__33368\,
            I => \N__33361\
        );

    \I__5852\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33358\
        );

    \I__5851\ : Span4Mux_v
    port map (
            O => \N__33364\,
            I => \N__33352\
        );

    \I__5850\ : Span4Mux_h
    port map (
            O => \N__33361\,
            I => \N__33352\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__33358\,
            I => \N__33349\
        );

    \I__5848\ : InMux
    port map (
            O => \N__33357\,
            I => \N__33346\
        );

    \I__5847\ : Span4Mux_v
    port map (
            O => \N__33352\,
            I => \N__33343\
        );

    \I__5846\ : Span4Mux_v
    port map (
            O => \N__33349\,
            I => \N__33338\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__33346\,
            I => \N__33338\
        );

    \I__5844\ : Odrv4
    port map (
            O => \N__33343\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__5843\ : Odrv4
    port map (
            O => \N__33338\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__5842\ : InMux
    port map (
            O => \N__33333\,
            I => \N__33329\
        );

    \I__5841\ : CascadeMux
    port map (
            O => \N__33332\,
            I => \N__33325\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__33329\,
            I => \N__33322\
        );

    \I__5839\ : InMux
    port map (
            O => \N__33328\,
            I => \N__33319\
        );

    \I__5838\ : InMux
    port map (
            O => \N__33325\,
            I => \N__33316\
        );

    \I__5837\ : Span4Mux_v
    port map (
            O => \N__33322\,
            I => \N__33313\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__33319\,
            I => \N__33310\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__33316\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__5834\ : Odrv4
    port map (
            O => \N__33313\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__5833\ : Odrv4
    port map (
            O => \N__33310\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__5832\ : CascadeMux
    port map (
            O => \N__33303\,
            I => \N__33300\
        );

    \I__5831\ : InMux
    port map (
            O => \N__33300\,
            I => \N__33297\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__33297\,
            I => \N__33294\
        );

    \I__5829\ : Span4Mux_v
    port map (
            O => \N__33294\,
            I => \N__33291\
        );

    \I__5828\ : Span4Mux_h
    port map (
            O => \N__33291\,
            I => \N__33288\
        );

    \I__5827\ : Odrv4
    port map (
            O => \N__33288\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\
        );

    \I__5826\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33282\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__33282\,
            I => \N__33277\
        );

    \I__5824\ : CascadeMux
    port map (
            O => \N__33281\,
            I => \N__33274\
        );

    \I__5823\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33271\
        );

    \I__5822\ : Span4Mux_h
    port map (
            O => \N__33277\,
            I => \N__33268\
        );

    \I__5821\ : InMux
    port map (
            O => \N__33274\,
            I => \N__33265\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__33271\,
            I => \N__33262\
        );

    \I__5819\ : Odrv4
    port map (
            O => \N__33268\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__33265\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__5817\ : Odrv4
    port map (
            O => \N__33262\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__5816\ : CascadeMux
    port map (
            O => \N__33255\,
            I => \N__33252\
        );

    \I__5815\ : InMux
    port map (
            O => \N__33252\,
            I => \N__33249\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__33249\,
            I => \N__33245\
        );

    \I__5813\ : InMux
    port map (
            O => \N__33248\,
            I => \N__33242\
        );

    \I__5812\ : Span4Mux_h
    port map (
            O => \N__33245\,
            I => \N__33238\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__33242\,
            I => \N__33235\
        );

    \I__5810\ : InMux
    port map (
            O => \N__33241\,
            I => \N__33232\
        );

    \I__5809\ : Span4Mux_v
    port map (
            O => \N__33238\,
            I => \N__33226\
        );

    \I__5808\ : Span4Mux_h
    port map (
            O => \N__33235\,
            I => \N__33226\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__33232\,
            I => \N__33223\
        );

    \I__5806\ : InMux
    port map (
            O => \N__33231\,
            I => \N__33220\
        );

    \I__5805\ : Span4Mux_v
    port map (
            O => \N__33226\,
            I => \N__33217\
        );

    \I__5804\ : Sp12to4
    port map (
            O => \N__33223\,
            I => \N__33212\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__33220\,
            I => \N__33212\
        );

    \I__5802\ : Odrv4
    port map (
            O => \N__33217\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__5801\ : Odrv12
    port map (
            O => \N__33212\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__5800\ : CascadeMux
    port map (
            O => \N__33207\,
            I => \N__33204\
        );

    \I__5799\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33201\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__33201\,
            I => \N__33198\
        );

    \I__5797\ : Span4Mux_v
    port map (
            O => \N__33198\,
            I => \N__33195\
        );

    \I__5796\ : Span4Mux_h
    port map (
            O => \N__33195\,
            I => \N__33192\
        );

    \I__5795\ : Odrv4
    port map (
            O => \N__33192\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\
        );

    \I__5794\ : InMux
    port map (
            O => \N__33189\,
            I => \N__33186\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__33186\,
            I => \N__33182\
        );

    \I__5792\ : CascadeMux
    port map (
            O => \N__33185\,
            I => \N__33178\
        );

    \I__5791\ : Span4Mux_h
    port map (
            O => \N__33182\,
            I => \N__33175\
        );

    \I__5790\ : InMux
    port map (
            O => \N__33181\,
            I => \N__33172\
        );

    \I__5789\ : InMux
    port map (
            O => \N__33178\,
            I => \N__33169\
        );

    \I__5788\ : Odrv4
    port map (
            O => \N__33175\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__33172\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__33169\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__5785\ : InMux
    port map (
            O => \N__33162\,
            I => \N__33158\
        );

    \I__5784\ : InMux
    port map (
            O => \N__33161\,
            I => \N__33155\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__33158\,
            I => \N__33151\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__33155\,
            I => \N__33148\
        );

    \I__5781\ : InMux
    port map (
            O => \N__33154\,
            I => \N__33145\
        );

    \I__5780\ : Span4Mux_v
    port map (
            O => \N__33151\,
            I => \N__33140\
        );

    \I__5779\ : Span4Mux_v
    port map (
            O => \N__33148\,
            I => \N__33140\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__33145\,
            I => \N__33137\
        );

    \I__5777\ : Span4Mux_h
    port map (
            O => \N__33140\,
            I => \N__33133\
        );

    \I__5776\ : Span4Mux_h
    port map (
            O => \N__33137\,
            I => \N__33130\
        );

    \I__5775\ : InMux
    port map (
            O => \N__33136\,
            I => \N__33127\
        );

    \I__5774\ : Odrv4
    port map (
            O => \N__33133\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__5773\ : Odrv4
    port map (
            O => \N__33130\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__33127\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__5771\ : CascadeMux
    port map (
            O => \N__33120\,
            I => \N__33117\
        );

    \I__5770\ : InMux
    port map (
            O => \N__33117\,
            I => \N__33114\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__33114\,
            I => \N__33111\
        );

    \I__5768\ : Span4Mux_v
    port map (
            O => \N__33111\,
            I => \N__33108\
        );

    \I__5767\ : Odrv4
    port map (
            O => \N__33108\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt26\
        );

    \I__5766\ : InMux
    port map (
            O => \N__33105\,
            I => \N__33101\
        );

    \I__5765\ : CascadeMux
    port map (
            O => \N__33104\,
            I => \N__33097\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__33101\,
            I => \N__33091\
        );

    \I__5763\ : InMux
    port map (
            O => \N__33100\,
            I => \N__33086\
        );

    \I__5762\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33086\
        );

    \I__5761\ : InMux
    port map (
            O => \N__33096\,
            I => \N__33083\
        );

    \I__5760\ : InMux
    port map (
            O => \N__33095\,
            I => \N__33078\
        );

    \I__5759\ : InMux
    port map (
            O => \N__33094\,
            I => \N__33078\
        );

    \I__5758\ : Span4Mux_h
    port map (
            O => \N__33091\,
            I => \N__33075\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__33086\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__33083\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__33078\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5754\ : Odrv4
    port map (
            O => \N__33075\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5753\ : InMux
    port map (
            O => \N__33066\,
            I => \N__33063\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__33063\,
            I => \N__33060\
        );

    \I__5751\ : Span4Mux_v
    port map (
            O => \N__33060\,
            I => \N__33057\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__33057\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_10\
        );

    \I__5749\ : InMux
    port map (
            O => \N__33054\,
            I => \N__33051\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__33051\,
            I => \N__33048\
        );

    \I__5747\ : Span4Mux_v
    port map (
            O => \N__33048\,
            I => \N__33045\
        );

    \I__5746\ : Odrv4
    port map (
            O => \N__33045\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_0\
        );

    \I__5745\ : InMux
    port map (
            O => \N__33042\,
            I => \N__33039\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__33039\,
            I => \N__33036\
        );

    \I__5743\ : Span4Mux_v
    port map (
            O => \N__33036\,
            I => \N__33033\
        );

    \I__5742\ : Odrv4
    port map (
            O => \N__33033\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_11\
        );

    \I__5741\ : CascadeMux
    port map (
            O => \N__33030\,
            I => \N__33026\
        );

    \I__5740\ : CascadeMux
    port map (
            O => \N__33029\,
            I => \N__33023\
        );

    \I__5739\ : InMux
    port map (
            O => \N__33026\,
            I => \N__33018\
        );

    \I__5738\ : InMux
    port map (
            O => \N__33023\,
            I => \N__33018\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__33018\,
            I => \N__33015\
        );

    \I__5736\ : Span4Mux_h
    port map (
            O => \N__33015\,
            I => \N__33012\
        );

    \I__5735\ : Odrv4
    port map (
            O => \N__33012\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_24\
        );

    \I__5734\ : InMux
    port map (
            O => \N__33009\,
            I => \N__33006\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__33006\,
            I => \N__33003\
        );

    \I__5732\ : Span4Mux_v
    port map (
            O => \N__33003\,
            I => \N__33000\
        );

    \I__5731\ : Span4Mux_h
    port map (
            O => \N__33000\,
            I => \N__32997\
        );

    \I__5730\ : Span4Mux_h
    port map (
            O => \N__32997\,
            I => \N__32994\
        );

    \I__5729\ : Odrv4
    port map (
            O => \N__32994\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_6\
        );

    \I__5728\ : InMux
    port map (
            O => \N__32991\,
            I => \N__32988\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__32988\,
            I => \N__32985\
        );

    \I__5726\ : Span4Mux_v
    port map (
            O => \N__32985\,
            I => \N__32982\
        );

    \I__5725\ : Odrv4
    port map (
            O => \N__32982\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_12\
        );

    \I__5724\ : InMux
    port map (
            O => \N__32979\,
            I => \N__32976\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__32976\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt22\
        );

    \I__5722\ : InMux
    port map (
            O => \N__32973\,
            I => \N__32968\
        );

    \I__5721\ : InMux
    port map (
            O => \N__32972\,
            I => \N__32963\
        );

    \I__5720\ : InMux
    port map (
            O => \N__32971\,
            I => \N__32963\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__32968\,
            I => \N__32958\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__32963\,
            I => \N__32958\
        );

    \I__5717\ : Odrv4
    port map (
            O => \N__32958\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_23\
        );

    \I__5716\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32950\
        );

    \I__5715\ : InMux
    port map (
            O => \N__32954\,
            I => \N__32945\
        );

    \I__5714\ : InMux
    port map (
            O => \N__32953\,
            I => \N__32945\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__32950\,
            I => \N__32940\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__32945\,
            I => \N__32940\
        );

    \I__5711\ : Odrv4
    port map (
            O => \N__32940\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_22\
        );

    \I__5710\ : CascadeMux
    port map (
            O => \N__32937\,
            I => \N__32934\
        );

    \I__5709\ : InMux
    port map (
            O => \N__32934\,
            I => \N__32931\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__32931\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22\
        );

    \I__5707\ : InMux
    port map (
            O => \N__32928\,
            I => \N__32925\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__32925\,
            I => \N__32922\
        );

    \I__5705\ : Span4Mux_h
    port map (
            O => \N__32922\,
            I => \N__32919\
        );

    \I__5704\ : Odrv4
    port map (
            O => \N__32919\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_4\
        );

    \I__5703\ : InMux
    port map (
            O => \N__32916\,
            I => \N__32913\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__32913\,
            I => \N__32910\
        );

    \I__5701\ : Odrv4
    port map (
            O => \N__32910\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_9\
        );

    \I__5700\ : InMux
    port map (
            O => \N__32907\,
            I => \N__32904\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__32904\,
            I => \N__32901\
        );

    \I__5698\ : Odrv4
    port map (
            O => \N__32901\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_13\
        );

    \I__5697\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32892\
        );

    \I__5696\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32892\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__32892\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_17\
        );

    \I__5694\ : InMux
    port map (
            O => \N__32889\,
            I => \N__32883\
        );

    \I__5693\ : InMux
    port map (
            O => \N__32888\,
            I => \N__32883\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__32883\,
            I => \N__32880\
        );

    \I__5691\ : Odrv4
    port map (
            O => \N__32880\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_25\
        );

    \I__5690\ : InMux
    port map (
            O => \N__32877\,
            I => \N__32873\
        );

    \I__5689\ : InMux
    port map (
            O => \N__32876\,
            I => \N__32869\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__32873\,
            I => \N__32866\
        );

    \I__5687\ : InMux
    port map (
            O => \N__32872\,
            I => \N__32863\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__32869\,
            I => \N__32860\
        );

    \I__5685\ : Span4Mux_v
    port map (
            O => \N__32866\,
            I => \N__32857\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__32863\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_27\
        );

    \I__5683\ : Odrv4
    port map (
            O => \N__32860\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_27\
        );

    \I__5682\ : Odrv4
    port map (
            O => \N__32857\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_27\
        );

    \I__5681\ : CascadeMux
    port map (
            O => \N__32850\,
            I => \N__32846\
        );

    \I__5680\ : CascadeMux
    port map (
            O => \N__32849\,
            I => \N__32843\
        );

    \I__5679\ : InMux
    port map (
            O => \N__32846\,
            I => \N__32839\
        );

    \I__5678\ : InMux
    port map (
            O => \N__32843\,
            I => \N__32836\
        );

    \I__5677\ : InMux
    port map (
            O => \N__32842\,
            I => \N__32833\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__32839\,
            I => \N__32830\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__32836\,
            I => \N__32827\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__32833\,
            I => \N__32822\
        );

    \I__5673\ : Span4Mux_v
    port map (
            O => \N__32830\,
            I => \N__32822\
        );

    \I__5672\ : Odrv4
    port map (
            O => \N__32827\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_26\
        );

    \I__5671\ : Odrv4
    port map (
            O => \N__32822\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_26\
        );

    \I__5670\ : InMux
    port map (
            O => \N__32817\,
            I => \N__32810\
        );

    \I__5669\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32810\
        );

    \I__5668\ : InMux
    port map (
            O => \N__32815\,
            I => \N__32807\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__32810\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__32807\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__5665\ : InMux
    port map (
            O => \N__32802\,
            I => \N__32794\
        );

    \I__5664\ : InMux
    port map (
            O => \N__32801\,
            I => \N__32789\
        );

    \I__5663\ : InMux
    port map (
            O => \N__32800\,
            I => \N__32789\
        );

    \I__5662\ : InMux
    port map (
            O => \N__32799\,
            I => \N__32784\
        );

    \I__5661\ : InMux
    port map (
            O => \N__32798\,
            I => \N__32784\
        );

    \I__5660\ : CascadeMux
    port map (
            O => \N__32797\,
            I => \N__32781\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__32794\,
            I => \N__32778\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__32789\,
            I => \N__32775\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__32784\,
            I => \N__32772\
        );

    \I__5656\ : InMux
    port map (
            O => \N__32781\,
            I => \N__32769\
        );

    \I__5655\ : Span4Mux_v
    port map (
            O => \N__32778\,
            I => \N__32766\
        );

    \I__5654\ : Span4Mux_v
    port map (
            O => \N__32775\,
            I => \N__32761\
        );

    \I__5653\ : Span4Mux_v
    port map (
            O => \N__32772\,
            I => \N__32761\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__32769\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5651\ : Odrv4
    port map (
            O => \N__32766\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5650\ : Odrv4
    port map (
            O => \N__32761\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5649\ : InMux
    port map (
            O => \N__32754\,
            I => \N__32751\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__32751\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_3\
        );

    \I__5647\ : InMux
    port map (
            O => \N__32748\,
            I => \N__32745\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__32745\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_5\
        );

    \I__5645\ : InMux
    port map (
            O => \N__32742\,
            I => \N__32739\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__32739\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_2\
        );

    \I__5643\ : InMux
    port map (
            O => \N__32736\,
            I => \N__32733\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__32733\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_1\
        );

    \I__5641\ : InMux
    port map (
            O => \N__32730\,
            I => \N__32727\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__32727\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_8\
        );

    \I__5639\ : CascadeMux
    port map (
            O => \N__32724\,
            I => \N__32721\
        );

    \I__5638\ : InMux
    port map (
            O => \N__32721\,
            I => \N__32718\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__32718\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt20\
        );

    \I__5636\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32708\
        );

    \I__5635\ : InMux
    port map (
            O => \N__32714\,
            I => \N__32708\
        );

    \I__5634\ : InMux
    port map (
            O => \N__32713\,
            I => \N__32705\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__32708\,
            I => \N__32702\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__32705\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_21\
        );

    \I__5631\ : Odrv4
    port map (
            O => \N__32702\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_21\
        );

    \I__5630\ : InMux
    port map (
            O => \N__32697\,
            I => \N__32690\
        );

    \I__5629\ : InMux
    port map (
            O => \N__32696\,
            I => \N__32690\
        );

    \I__5628\ : InMux
    port map (
            O => \N__32695\,
            I => \N__32687\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__32690\,
            I => \N__32684\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__32687\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_20\
        );

    \I__5625\ : Odrv4
    port map (
            O => \N__32684\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_20\
        );

    \I__5624\ : InMux
    port map (
            O => \N__32679\,
            I => \N__32676\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__32676\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20\
        );

    \I__5622\ : CascadeMux
    port map (
            O => \N__32673\,
            I => \N__32670\
        );

    \I__5621\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32667\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__32667\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22\
        );

    \I__5619\ : InMux
    port map (
            O => \N__32664\,
            I => \N__32661\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__32661\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt20\
        );

    \I__5617\ : InMux
    port map (
            O => \N__32658\,
            I => \N__32655\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__32655\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt22\
        );

    \I__5615\ : CascadeMux
    port map (
            O => \N__32652\,
            I => \N__32649\
        );

    \I__5614\ : InMux
    port map (
            O => \N__32649\,
            I => \N__32646\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__32646\,
            I => \N__32643\
        );

    \I__5612\ : Odrv4
    port map (
            O => \N__32643\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20\
        );

    \I__5611\ : CascadeMux
    port map (
            O => \N__32640\,
            I => \N__32637\
        );

    \I__5610\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32634\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__32634\,
            I => \N__32631\
        );

    \I__5608\ : Odrv4
    port map (
            O => \N__32631\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24\
        );

    \I__5607\ : InMux
    port map (
            O => \N__32628\,
            I => \N__32625\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__32625\,
            I => \N__32622\
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__32622\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt30\
        );

    \I__5604\ : InMux
    port map (
            O => \N__32619\,
            I => \N__32616\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__32616\,
            I => \N__32613\
        );

    \I__5602\ : Odrv4
    port map (
            O => \N__32613\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt24\
        );

    \I__5601\ : CEMux
    port map (
            O => \N__32610\,
            I => \N__32606\
        );

    \I__5600\ : CEMux
    port map (
            O => \N__32609\,
            I => \N__32603\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__32606\,
            I => \N__32599\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__32603\,
            I => \N__32595\
        );

    \I__5597\ : CEMux
    port map (
            O => \N__32602\,
            I => \N__32592\
        );

    \I__5596\ : Span4Mux_h
    port map (
            O => \N__32599\,
            I => \N__32589\
        );

    \I__5595\ : CEMux
    port map (
            O => \N__32598\,
            I => \N__32586\
        );

    \I__5594\ : Span4Mux_h
    port map (
            O => \N__32595\,
            I => \N__32583\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__32592\,
            I => \N__32580\
        );

    \I__5592\ : Span4Mux_v
    port map (
            O => \N__32589\,
            I => \N__32577\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__32586\,
            I => \N__32574\
        );

    \I__5590\ : Span4Mux_v
    port map (
            O => \N__32583\,
            I => \N__32571\
        );

    \I__5589\ : Span4Mux_h
    port map (
            O => \N__32580\,
            I => \N__32568\
        );

    \I__5588\ : Span4Mux_v
    port map (
            O => \N__32577\,
            I => \N__32565\
        );

    \I__5587\ : Span12Mux_v
    port map (
            O => \N__32574\,
            I => \N__32562\
        );

    \I__5586\ : Sp12to4
    port map (
            O => \N__32571\,
            I => \N__32557\
        );

    \I__5585\ : Sp12to4
    port map (
            O => \N__32568\,
            I => \N__32557\
        );

    \I__5584\ : Odrv4
    port map (
            O => \N__32565\,
            I => \current_shift_inst.timer_s1.N_154_i\
        );

    \I__5583\ : Odrv12
    port map (
            O => \N__32562\,
            I => \current_shift_inst.timer_s1.N_154_i\
        );

    \I__5582\ : Odrv12
    port map (
            O => \N__32557\,
            I => \current_shift_inst.timer_s1.N_154_i\
        );

    \I__5581\ : CascadeMux
    port map (
            O => \N__32550\,
            I => \N__32547\
        );

    \I__5580\ : InMux
    port map (
            O => \N__32547\,
            I => \N__32544\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__32544\,
            I => \N__32541\
        );

    \I__5578\ : Span4Mux_v
    port map (
            O => \N__32541\,
            I => \N__32538\
        );

    \I__5577\ : Odrv4
    port map (
            O => \N__32538\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30\
        );

    \I__5576\ : CascadeMux
    port map (
            O => \N__32535\,
            I => \N__32532\
        );

    \I__5575\ : InMux
    port map (
            O => \N__32532\,
            I => \N__32529\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__32529\,
            I => \N__32526\
        );

    \I__5573\ : Odrv12
    port map (
            O => \N__32526\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt26\
        );

    \I__5572\ : InMux
    port map (
            O => \N__32523\,
            I => \N__32520\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__32520\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28\
        );

    \I__5570\ : InMux
    port map (
            O => \N__32517\,
            I => \bfn_11_28_0_\
        );

    \I__5569\ : CascadeMux
    port map (
            O => \N__32514\,
            I => \N__32511\
        );

    \I__5568\ : InMux
    port map (
            O => \N__32511\,
            I => \N__32508\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__32508\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt28\
        );

    \I__5566\ : CascadeMux
    port map (
            O => \N__32505\,
            I => \N__32502\
        );

    \I__5565\ : InMux
    port map (
            O => \N__32502\,
            I => \N__32499\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__32499\,
            I => \phase_controller_inst1.stoper_tr.counter_i_10\
        );

    \I__5563\ : CascadeMux
    port map (
            O => \N__32496\,
            I => \N__32493\
        );

    \I__5562\ : InMux
    port map (
            O => \N__32493\,
            I => \N__32490\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__32490\,
            I => \N__32487\
        );

    \I__5560\ : Odrv4
    port map (
            O => \N__32487\,
            I => \phase_controller_inst1.stoper_tr.counter_i_11\
        );

    \I__5559\ : CascadeMux
    port map (
            O => \N__32484\,
            I => \N__32481\
        );

    \I__5558\ : InMux
    port map (
            O => \N__32481\,
            I => \N__32478\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__32478\,
            I => \N__32475\
        );

    \I__5556\ : Odrv4
    port map (
            O => \N__32475\,
            I => \phase_controller_inst1.stoper_tr.counter_i_12\
        );

    \I__5555\ : CascadeMux
    port map (
            O => \N__32472\,
            I => \N__32469\
        );

    \I__5554\ : InMux
    port map (
            O => \N__32469\,
            I => \N__32466\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__32466\,
            I => \N__32463\
        );

    \I__5552\ : Odrv4
    port map (
            O => \N__32463\,
            I => \phase_controller_inst1.stoper_tr.counter_i_13\
        );

    \I__5551\ : CascadeMux
    port map (
            O => \N__32460\,
            I => \N__32457\
        );

    \I__5550\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32454\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__32454\,
            I => \N__32451\
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__32451\,
            I => \phase_controller_inst1.stoper_tr.counter_i_14\
        );

    \I__5547\ : CascadeMux
    port map (
            O => \N__32448\,
            I => \N__32445\
        );

    \I__5546\ : InMux
    port map (
            O => \N__32445\,
            I => \N__32442\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__32442\,
            I => \phase_controller_inst1.stoper_tr.counter_i_15\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__32439\,
            I => \N__32436\
        );

    \I__5543\ : InMux
    port map (
            O => \N__32436\,
            I => \N__32433\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__32433\,
            I => \phase_controller_inst1.stoper_tr.counter_i_1\
        );

    \I__5541\ : CascadeMux
    port map (
            O => \N__32430\,
            I => \N__32427\
        );

    \I__5540\ : InMux
    port map (
            O => \N__32427\,
            I => \N__32424\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__32424\,
            I => \phase_controller_inst1.stoper_tr.counter_i_2\
        );

    \I__5538\ : CascadeMux
    port map (
            O => \N__32421\,
            I => \N__32418\
        );

    \I__5537\ : InMux
    port map (
            O => \N__32418\,
            I => \N__32415\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__32415\,
            I => \phase_controller_inst1.stoper_tr.counter_i_3\
        );

    \I__5535\ : CascadeMux
    port map (
            O => \N__32412\,
            I => \N__32409\
        );

    \I__5534\ : InMux
    port map (
            O => \N__32409\,
            I => \N__32406\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__32406\,
            I => \N__32403\
        );

    \I__5532\ : Odrv4
    port map (
            O => \N__32403\,
            I => \phase_controller_inst1.stoper_tr.counter_i_4\
        );

    \I__5531\ : CascadeMux
    port map (
            O => \N__32400\,
            I => \N__32397\
        );

    \I__5530\ : InMux
    port map (
            O => \N__32397\,
            I => \N__32394\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__32394\,
            I => \phase_controller_inst1.stoper_tr.counter_i_5\
        );

    \I__5528\ : CascadeMux
    port map (
            O => \N__32391\,
            I => \N__32388\
        );

    \I__5527\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32385\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__32385\,
            I => \N__32382\
        );

    \I__5525\ : Odrv4
    port map (
            O => \N__32382\,
            I => \phase_controller_inst1.stoper_tr.counter_i_6\
        );

    \I__5524\ : CascadeMux
    port map (
            O => \N__32379\,
            I => \N__32376\
        );

    \I__5523\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32373\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__32373\,
            I => \phase_controller_inst1.stoper_tr.counter_i_7\
        );

    \I__5521\ : CascadeMux
    port map (
            O => \N__32370\,
            I => \N__32367\
        );

    \I__5520\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32364\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__32364\,
            I => \phase_controller_inst1.stoper_tr.counter_i_8\
        );

    \I__5518\ : CascadeMux
    port map (
            O => \N__32361\,
            I => \N__32358\
        );

    \I__5517\ : InMux
    port map (
            O => \N__32358\,
            I => \N__32355\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__32355\,
            I => \phase_controller_inst1.stoper_tr.counter_i_9\
        );

    \I__5515\ : CascadeMux
    port map (
            O => \N__32352\,
            I => \N__32349\
        );

    \I__5514\ : InMux
    port map (
            O => \N__32349\,
            I => \N__32346\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__32346\,
            I => \N__32342\
        );

    \I__5512\ : InMux
    port map (
            O => \N__32345\,
            I => \N__32339\
        );

    \I__5511\ : Span4Mux_h
    port map (
            O => \N__32342\,
            I => \N__32335\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__32339\,
            I => \N__32332\
        );

    \I__5509\ : InMux
    port map (
            O => \N__32338\,
            I => \N__32329\
        );

    \I__5508\ : Span4Mux_v
    port map (
            O => \N__32335\,
            I => \N__32323\
        );

    \I__5507\ : Span4Mux_h
    port map (
            O => \N__32332\,
            I => \N__32323\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__32329\,
            I => \N__32320\
        );

    \I__5505\ : InMux
    port map (
            O => \N__32328\,
            I => \N__32317\
        );

    \I__5504\ : Odrv4
    port map (
            O => \N__32323\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__5503\ : Odrv12
    port map (
            O => \N__32320\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__32317\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__5501\ : InMux
    port map (
            O => \N__32310\,
            I => \N__32307\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__32307\,
            I => \N__32304\
        );

    \I__5499\ : Odrv12
    port map (
            O => \N__32304\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__5498\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32297\
        );

    \I__5497\ : CascadeMux
    port map (
            O => \N__32300\,
            I => \N__32294\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__32297\,
            I => \N__32290\
        );

    \I__5495\ : InMux
    port map (
            O => \N__32294\,
            I => \N__32287\
        );

    \I__5494\ : InMux
    port map (
            O => \N__32293\,
            I => \N__32284\
        );

    \I__5493\ : Span4Mux_v
    port map (
            O => \N__32290\,
            I => \N__32277\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__32287\,
            I => \N__32277\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__32284\,
            I => \N__32277\
        );

    \I__5490\ : Span4Mux_v
    port map (
            O => \N__32277\,
            I => \N__32273\
        );

    \I__5489\ : InMux
    port map (
            O => \N__32276\,
            I => \N__32270\
        );

    \I__5488\ : Odrv4
    port map (
            O => \N__32273\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__32270\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__5486\ : InMux
    port map (
            O => \N__32265\,
            I => \N__32262\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__32262\,
            I => \N__32259\
        );

    \I__5484\ : Odrv12
    port map (
            O => \N__32259\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__5483\ : InMux
    port map (
            O => \N__32256\,
            I => \N__32253\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__32253\,
            I => \N__32248\
        );

    \I__5481\ : InMux
    port map (
            O => \N__32252\,
            I => \N__32245\
        );

    \I__5480\ : InMux
    port map (
            O => \N__32251\,
            I => \N__32242\
        );

    \I__5479\ : Span4Mux_v
    port map (
            O => \N__32248\,
            I => \N__32235\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__32245\,
            I => \N__32235\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__32242\,
            I => \N__32235\
        );

    \I__5476\ : Span4Mux_v
    port map (
            O => \N__32235\,
            I => \N__32231\
        );

    \I__5475\ : InMux
    port map (
            O => \N__32234\,
            I => \N__32228\
        );

    \I__5474\ : Odrv4
    port map (
            O => \N__32231\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__32228\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__5472\ : InMux
    port map (
            O => \N__32223\,
            I => \N__32220\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__32220\,
            I => \N__32217\
        );

    \I__5470\ : Span4Mux_v
    port map (
            O => \N__32217\,
            I => \N__32214\
        );

    \I__5469\ : Odrv4
    port map (
            O => \N__32214\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__5468\ : CascadeMux
    port map (
            O => \N__32211\,
            I => \N__32208\
        );

    \I__5467\ : InMux
    port map (
            O => \N__32208\,
            I => \N__32205\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__32205\,
            I => \N__32201\
        );

    \I__5465\ : InMux
    port map (
            O => \N__32204\,
            I => \N__32198\
        );

    \I__5464\ : Span4Mux_v
    port map (
            O => \N__32201\,
            I => \N__32192\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__32198\,
            I => \N__32192\
        );

    \I__5462\ : InMux
    port map (
            O => \N__32197\,
            I => \N__32189\
        );

    \I__5461\ : Span4Mux_h
    port map (
            O => \N__32192\,
            I => \N__32186\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__32189\,
            I => \N__32183\
        );

    \I__5459\ : Span4Mux_v
    port map (
            O => \N__32186\,
            I => \N__32179\
        );

    \I__5458\ : Span4Mux_v
    port map (
            O => \N__32183\,
            I => \N__32176\
        );

    \I__5457\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32173\
        );

    \I__5456\ : Odrv4
    port map (
            O => \N__32179\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__5455\ : Odrv4
    port map (
            O => \N__32176\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__32173\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__5453\ : InMux
    port map (
            O => \N__32166\,
            I => \N__32163\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__32163\,
            I => \N__32160\
        );

    \I__5451\ : Odrv12
    port map (
            O => \N__32160\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__32157\,
            I => \N__32154\
        );

    \I__5449\ : InMux
    port map (
            O => \N__32154\,
            I => \N__32151\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__32151\,
            I => \N__32146\
        );

    \I__5447\ : InMux
    port map (
            O => \N__32150\,
            I => \N__32141\
        );

    \I__5446\ : InMux
    port map (
            O => \N__32149\,
            I => \N__32141\
        );

    \I__5445\ : Span4Mux_v
    port map (
            O => \N__32146\,
            I => \N__32135\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__32141\,
            I => \N__32135\
        );

    \I__5443\ : InMux
    port map (
            O => \N__32140\,
            I => \N__32132\
        );

    \I__5442\ : Span4Mux_v
    port map (
            O => \N__32135\,
            I => \N__32129\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__32132\,
            I => \N__32126\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__32129\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__5439\ : Odrv4
    port map (
            O => \N__32126\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__5438\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32118\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__32118\,
            I => \N__32115\
        );

    \I__5436\ : Span4Mux_v
    port map (
            O => \N__32115\,
            I => \N__32112\
        );

    \I__5435\ : Span4Mux_v
    port map (
            O => \N__32112\,
            I => \N__32109\
        );

    \I__5434\ : Odrv4
    port map (
            O => \N__32109\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__5433\ : InMux
    port map (
            O => \N__32106\,
            I => \N__32103\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__32103\,
            I => \N__32099\
        );

    \I__5431\ : InMux
    port map (
            O => \N__32102\,
            I => \N__32095\
        );

    \I__5430\ : Span4Mux_h
    port map (
            O => \N__32099\,
            I => \N__32092\
        );

    \I__5429\ : InMux
    port map (
            O => \N__32098\,
            I => \N__32089\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__32095\,
            I => \N__32085\
        );

    \I__5427\ : Span4Mux_v
    port map (
            O => \N__32092\,
            I => \N__32080\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__32089\,
            I => \N__32080\
        );

    \I__5425\ : InMux
    port map (
            O => \N__32088\,
            I => \N__32077\
        );

    \I__5424\ : Span4Mux_v
    port map (
            O => \N__32085\,
            I => \N__32074\
        );

    \I__5423\ : Span4Mux_v
    port map (
            O => \N__32080\,
            I => \N__32069\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__32077\,
            I => \N__32069\
        );

    \I__5421\ : Odrv4
    port map (
            O => \N__32074\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__5420\ : Odrv4
    port map (
            O => \N__32069\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__5419\ : InMux
    port map (
            O => \N__32064\,
            I => \N__32061\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__32061\,
            I => \N__32058\
        );

    \I__5417\ : Sp12to4
    port map (
            O => \N__32058\,
            I => \N__32055\
        );

    \I__5416\ : Odrv12
    port map (
            O => \N__32055\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__5415\ : InMux
    port map (
            O => \N__32052\,
            I => \N__32049\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__32049\,
            I => \phase_controller_inst1.stoper_tr.counter_i_0\
        );

    \I__5413\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32043\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__32043\,
            I => \N__32040\
        );

    \I__5411\ : Span4Mux_h
    port map (
            O => \N__32040\,
            I => \N__32037\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__32037\,
            I => \N__32034\
        );

    \I__5409\ : Span4Mux_v
    port map (
            O => \N__32034\,
            I => \N__32031\
        );

    \I__5408\ : Odrv4
    port map (
            O => \N__32031\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__5407\ : CascadeMux
    port map (
            O => \N__32028\,
            I => \N__32025\
        );

    \I__5406\ : InMux
    port map (
            O => \N__32025\,
            I => \N__32022\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__32022\,
            I => \N__32019\
        );

    \I__5404\ : Span4Mux_h
    port map (
            O => \N__32019\,
            I => \N__32013\
        );

    \I__5403\ : InMux
    port map (
            O => \N__32018\,
            I => \N__32008\
        );

    \I__5402\ : InMux
    port map (
            O => \N__32017\,
            I => \N__32008\
        );

    \I__5401\ : InMux
    port map (
            O => \N__32016\,
            I => \N__32005\
        );

    \I__5400\ : Sp12to4
    port map (
            O => \N__32013\,
            I => \N__32002\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__32008\,
            I => \N__31999\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__32005\,
            I => \N__31996\
        );

    \I__5397\ : Span12Mux_v
    port map (
            O => \N__32002\,
            I => \N__31993\
        );

    \I__5396\ : Span4Mux_h
    port map (
            O => \N__31999\,
            I => \N__31990\
        );

    \I__5395\ : Odrv4
    port map (
            O => \N__31996\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__5394\ : Odrv12
    port map (
            O => \N__31993\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__5393\ : Odrv4
    port map (
            O => \N__31990\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__5392\ : InMux
    port map (
            O => \N__31983\,
            I => \bfn_11_22_0_\
        );

    \I__5391\ : InMux
    port map (
            O => \N__31980\,
            I => \N__31977\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__31977\,
            I => \N__31974\
        );

    \I__5389\ : Span4Mux_h
    port map (
            O => \N__31974\,
            I => \N__31971\
        );

    \I__5388\ : Span4Mux_h
    port map (
            O => \N__31971\,
            I => \N__31968\
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__31968\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\
        );

    \I__5386\ : CascadeMux
    port map (
            O => \N__31965\,
            I => \N__31962\
        );

    \I__5385\ : InMux
    port map (
            O => \N__31962\,
            I => \N__31959\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__31959\,
            I => \N__31955\
        );

    \I__5383\ : CascadeMux
    port map (
            O => \N__31958\,
            I => \N__31950\
        );

    \I__5382\ : Span4Mux_v
    port map (
            O => \N__31955\,
            I => \N__31947\
        );

    \I__5381\ : InMux
    port map (
            O => \N__31954\,
            I => \N__31944\
        );

    \I__5380\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31939\
        );

    \I__5379\ : InMux
    port map (
            O => \N__31950\,
            I => \N__31939\
        );

    \I__5378\ : Span4Mux_v
    port map (
            O => \N__31947\,
            I => \N__31936\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__31944\,
            I => \N__31931\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__31939\,
            I => \N__31931\
        );

    \I__5375\ : Sp12to4
    port map (
            O => \N__31936\,
            I => \N__31928\
        );

    \I__5374\ : Span4Mux_h
    port map (
            O => \N__31931\,
            I => \N__31925\
        );

    \I__5373\ : Odrv12
    port map (
            O => \N__31928\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__5372\ : Odrv4
    port map (
            O => \N__31925\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__5371\ : InMux
    port map (
            O => \N__31920\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__5370\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31914\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__31914\,
            I => \N__31911\
        );

    \I__5368\ : Span4Mux_h
    port map (
            O => \N__31911\,
            I => \N__31908\
        );

    \I__5367\ : Span4Mux_h
    port map (
            O => \N__31908\,
            I => \N__31905\
        );

    \I__5366\ : Span4Mux_v
    port map (
            O => \N__31905\,
            I => \N__31902\
        );

    \I__5365\ : Odrv4
    port map (
            O => \N__31902\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\
        );

    \I__5364\ : CascadeMux
    port map (
            O => \N__31899\,
            I => \N__31896\
        );

    \I__5363\ : InMux
    port map (
            O => \N__31896\,
            I => \N__31893\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__31893\,
            I => \N__31890\
        );

    \I__5361\ : Span4Mux_h
    port map (
            O => \N__31890\,
            I => \N__31887\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__31887\,
            I => \N__31883\
        );

    \I__5359\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31879\
        );

    \I__5358\ : Sp12to4
    port map (
            O => \N__31883\,
            I => \N__31875\
        );

    \I__5357\ : InMux
    port map (
            O => \N__31882\,
            I => \N__31872\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__31879\,
            I => \N__31869\
        );

    \I__5355\ : InMux
    port map (
            O => \N__31878\,
            I => \N__31866\
        );

    \I__5354\ : Span12Mux_v
    port map (
            O => \N__31875\,
            I => \N__31863\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__31872\,
            I => \N__31858\
        );

    \I__5352\ : Span4Mux_v
    port map (
            O => \N__31869\,
            I => \N__31858\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__31866\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5350\ : Odrv12
    port map (
            O => \N__31863\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5349\ : Odrv4
    port map (
            O => \N__31858\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5348\ : InMux
    port map (
            O => \N__31851\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__5347\ : InMux
    port map (
            O => \N__31848\,
            I => \N__31845\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__31845\,
            I => \N__31842\
        );

    \I__5345\ : Odrv12
    port map (
            O => \N__31842\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\
        );

    \I__5344\ : CascadeMux
    port map (
            O => \N__31839\,
            I => \N__31836\
        );

    \I__5343\ : InMux
    port map (
            O => \N__31836\,
            I => \N__31833\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__31833\,
            I => \N__31830\
        );

    \I__5341\ : Span4Mux_h
    port map (
            O => \N__31830\,
            I => \N__31827\
        );

    \I__5340\ : Span4Mux_h
    port map (
            O => \N__31827\,
            I => \N__31821\
        );

    \I__5339\ : CascadeMux
    port map (
            O => \N__31826\,
            I => \N__31818\
        );

    \I__5338\ : InMux
    port map (
            O => \N__31825\,
            I => \N__31815\
        );

    \I__5337\ : CascadeMux
    port map (
            O => \N__31824\,
            I => \N__31812\
        );

    \I__5336\ : Span4Mux_v
    port map (
            O => \N__31821\,
            I => \N__31809\
        );

    \I__5335\ : InMux
    port map (
            O => \N__31818\,
            I => \N__31806\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__31815\,
            I => \N__31803\
        );

    \I__5333\ : InMux
    port map (
            O => \N__31812\,
            I => \N__31800\
        );

    \I__5332\ : Span4Mux_v
    port map (
            O => \N__31809\,
            I => \N__31795\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__31806\,
            I => \N__31795\
        );

    \I__5330\ : Span4Mux_v
    port map (
            O => \N__31803\,
            I => \N__31792\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__31800\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__5328\ : Odrv4
    port map (
            O => \N__31795\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__5327\ : Odrv4
    port map (
            O => \N__31792\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__5326\ : InMux
    port map (
            O => \N__31785\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__5325\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31779\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__31779\,
            I => \N__31776\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__31776\,
            I => \N__31773\
        );

    \I__5322\ : Span4Mux_h
    port map (
            O => \N__31773\,
            I => \N__31770\
        );

    \I__5321\ : Span4Mux_v
    port map (
            O => \N__31770\,
            I => \N__31767\
        );

    \I__5320\ : Odrv4
    port map (
            O => \N__31767\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\
        );

    \I__5319\ : CascadeMux
    port map (
            O => \N__31764\,
            I => \N__31761\
        );

    \I__5318\ : InMux
    port map (
            O => \N__31761\,
            I => \N__31758\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__31758\,
            I => \N__31753\
        );

    \I__5316\ : InMux
    port map (
            O => \N__31757\,
            I => \N__31748\
        );

    \I__5315\ : InMux
    port map (
            O => \N__31756\,
            I => \N__31748\
        );

    \I__5314\ : Sp12to4
    port map (
            O => \N__31753\,
            I => \N__31744\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__31748\,
            I => \N__31741\
        );

    \I__5312\ : InMux
    port map (
            O => \N__31747\,
            I => \N__31738\
        );

    \I__5311\ : Span12Mux_v
    port map (
            O => \N__31744\,
            I => \N__31735\
        );

    \I__5310\ : Span4Mux_h
    port map (
            O => \N__31741\,
            I => \N__31732\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__31738\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__5308\ : Odrv12
    port map (
            O => \N__31735\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__5307\ : Odrv4
    port map (
            O => \N__31732\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__5306\ : InMux
    port map (
            O => \N__31725\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__5305\ : InMux
    port map (
            O => \N__31722\,
            I => \N__31719\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__31719\,
            I => \N__31716\
        );

    \I__5303\ : Odrv12
    port map (
            O => \N__31716\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\
        );

    \I__5302\ : CascadeMux
    port map (
            O => \N__31713\,
            I => \N__31710\
        );

    \I__5301\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31707\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__31707\,
            I => \N__31703\
        );

    \I__5299\ : CascadeMux
    port map (
            O => \N__31706\,
            I => \N__31700\
        );

    \I__5298\ : Span4Mux_h
    port map (
            O => \N__31703\,
            I => \N__31697\
        );

    \I__5297\ : InMux
    port map (
            O => \N__31700\,
            I => \N__31694\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__31697\,
            I => \N__31691\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__31694\,
            I => \N__31686\
        );

    \I__5294\ : Span4Mux_v
    port map (
            O => \N__31691\,
            I => \N__31683\
        );

    \I__5293\ : InMux
    port map (
            O => \N__31690\,
            I => \N__31680\
        );

    \I__5292\ : InMux
    port map (
            O => \N__31689\,
            I => \N__31677\
        );

    \I__5291\ : Span4Mux_h
    port map (
            O => \N__31686\,
            I => \N__31674\
        );

    \I__5290\ : Span4Mux_v
    port map (
            O => \N__31683\,
            I => \N__31669\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__31680\,
            I => \N__31669\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__31677\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__5287\ : Odrv4
    port map (
            O => \N__31674\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__5286\ : Odrv4
    port map (
            O => \N__31669\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__5285\ : InMux
    port map (
            O => \N__31662\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__5284\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31656\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__31656\,
            I => \N__31644\
        );

    \I__5282\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31637\
        );

    \I__5281\ : InMux
    port map (
            O => \N__31654\,
            I => \N__31626\
        );

    \I__5280\ : InMux
    port map (
            O => \N__31653\,
            I => \N__31626\
        );

    \I__5279\ : InMux
    port map (
            O => \N__31652\,
            I => \N__31626\
        );

    \I__5278\ : InMux
    port map (
            O => \N__31651\,
            I => \N__31626\
        );

    \I__5277\ : InMux
    port map (
            O => \N__31650\,
            I => \N__31617\
        );

    \I__5276\ : InMux
    port map (
            O => \N__31649\,
            I => \N__31617\
        );

    \I__5275\ : InMux
    port map (
            O => \N__31648\,
            I => \N__31617\
        );

    \I__5274\ : InMux
    port map (
            O => \N__31647\,
            I => \N__31617\
        );

    \I__5273\ : Span4Mux_v
    port map (
            O => \N__31644\,
            I => \N__31614\
        );

    \I__5272\ : InMux
    port map (
            O => \N__31643\,
            I => \N__31610\
        );

    \I__5271\ : InMux
    port map (
            O => \N__31642\,
            I => \N__31605\
        );

    \I__5270\ : InMux
    port map (
            O => \N__31641\,
            I => \N__31605\
        );

    \I__5269\ : InMux
    port map (
            O => \N__31640\,
            I => \N__31602\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__31637\,
            I => \N__31599\
        );

    \I__5267\ : InMux
    port map (
            O => \N__31636\,
            I => \N__31596\
        );

    \I__5266\ : InMux
    port map (
            O => \N__31635\,
            I => \N__31579\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__31626\,
            I => \N__31574\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__31617\,
            I => \N__31574\
        );

    \I__5263\ : Sp12to4
    port map (
            O => \N__31614\,
            I => \N__31571\
        );

    \I__5262\ : InMux
    port map (
            O => \N__31613\,
            I => \N__31568\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__31610\,
            I => \N__31563\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__31605\,
            I => \N__31563\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__31602\,
            I => \N__31560\
        );

    \I__5258\ : Span4Mux_v
    port map (
            O => \N__31599\,
            I => \N__31555\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__31596\,
            I => \N__31555\
        );

    \I__5256\ : InMux
    port map (
            O => \N__31595\,
            I => \N__31552\
        );

    \I__5255\ : InMux
    port map (
            O => \N__31594\,
            I => \N__31545\
        );

    \I__5254\ : InMux
    port map (
            O => \N__31593\,
            I => \N__31545\
        );

    \I__5253\ : InMux
    port map (
            O => \N__31592\,
            I => \N__31545\
        );

    \I__5252\ : InMux
    port map (
            O => \N__31591\,
            I => \N__31542\
        );

    \I__5251\ : InMux
    port map (
            O => \N__31590\,
            I => \N__31535\
        );

    \I__5250\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31535\
        );

    \I__5249\ : InMux
    port map (
            O => \N__31588\,
            I => \N__31535\
        );

    \I__5248\ : InMux
    port map (
            O => \N__31587\,
            I => \N__31522\
        );

    \I__5247\ : InMux
    port map (
            O => \N__31586\,
            I => \N__31522\
        );

    \I__5246\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31522\
        );

    \I__5245\ : InMux
    port map (
            O => \N__31584\,
            I => \N__31522\
        );

    \I__5244\ : InMux
    port map (
            O => \N__31583\,
            I => \N__31522\
        );

    \I__5243\ : InMux
    port map (
            O => \N__31582\,
            I => \N__31522\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__31579\,
            I => \N__31517\
        );

    \I__5241\ : Span4Mux_v
    port map (
            O => \N__31574\,
            I => \N__31517\
        );

    \I__5240\ : Span12Mux_h
    port map (
            O => \N__31571\,
            I => \N__31514\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__31568\,
            I => \N__31505\
        );

    \I__5238\ : Span4Mux_v
    port map (
            O => \N__31563\,
            I => \N__31505\
        );

    \I__5237\ : Span4Mux_h
    port map (
            O => \N__31560\,
            I => \N__31505\
        );

    \I__5236\ : Span4Mux_h
    port map (
            O => \N__31555\,
            I => \N__31505\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__31552\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__31545\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__31542\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__31535\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__31522\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5230\ : Odrv4
    port map (
            O => \N__31517\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5229\ : Odrv12
    port map (
            O => \N__31514\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5228\ : Odrv4
    port map (
            O => \N__31505\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5227\ : InMux
    port map (
            O => \N__31488\,
            I => \N__31485\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__31485\,
            I => \N__31482\
        );

    \I__5225\ : Span4Mux_h
    port map (
            O => \N__31482\,
            I => \N__31479\
        );

    \I__5224\ : Span4Mux_h
    port map (
            O => \N__31479\,
            I => \N__31476\
        );

    \I__5223\ : Odrv4
    port map (
            O => \N__31476\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\
        );

    \I__5222\ : InMux
    port map (
            O => \N__31473\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__5221\ : IoInMux
    port map (
            O => \N__31470\,
            I => \N__31467\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__31467\,
            I => \N__31464\
        );

    \I__5219\ : Span4Mux_s3_v
    port map (
            O => \N__31464\,
            I => \N__31461\
        );

    \I__5218\ : Span4Mux_h
    port map (
            O => \N__31461\,
            I => \N__31458\
        );

    \I__5217\ : Span4Mux_v
    port map (
            O => \N__31458\,
            I => \N__31455\
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__31455\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__5215\ : InMux
    port map (
            O => \N__31452\,
            I => \N__31449\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__31449\,
            I => \N__31446\
        );

    \I__5213\ : Odrv12
    port map (
            O => \N__31446\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__31443\,
            I => \N__31440\
        );

    \I__5211\ : InMux
    port map (
            O => \N__31440\,
            I => \N__31437\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__31437\,
            I => \N__31433\
        );

    \I__5209\ : CascadeMux
    port map (
            O => \N__31436\,
            I => \N__31430\
        );

    \I__5208\ : Span4Mux_v
    port map (
            O => \N__31433\,
            I => \N__31426\
        );

    \I__5207\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31423\
        );

    \I__5206\ : InMux
    port map (
            O => \N__31429\,
            I => \N__31420\
        );

    \I__5205\ : Sp12to4
    port map (
            O => \N__31426\,
            I => \N__31416\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__31423\,
            I => \N__31413\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__31420\,
            I => \N__31410\
        );

    \I__5202\ : InMux
    port map (
            O => \N__31419\,
            I => \N__31407\
        );

    \I__5201\ : Span12Mux_h
    port map (
            O => \N__31416\,
            I => \N__31404\
        );

    \I__5200\ : Span4Mux_h
    port map (
            O => \N__31413\,
            I => \N__31399\
        );

    \I__5199\ : Span4Mux_h
    port map (
            O => \N__31410\,
            I => \N__31399\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__31407\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5197\ : Odrv12
    port map (
            O => \N__31404\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5196\ : Odrv4
    port map (
            O => \N__31399\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5195\ : InMux
    port map (
            O => \N__31392\,
            I => \bfn_11_21_0_\
        );

    \I__5194\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31386\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__31386\,
            I => \N__31383\
        );

    \I__5192\ : Span4Mux_h
    port map (
            O => \N__31383\,
            I => \N__31380\
        );

    \I__5191\ : Span4Mux_h
    port map (
            O => \N__31380\,
            I => \N__31377\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__31377\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__31374\,
            I => \N__31371\
        );

    \I__5188\ : InMux
    port map (
            O => \N__31371\,
            I => \N__31368\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__31368\,
            I => \N__31365\
        );

    \I__5186\ : Span4Mux_h
    port map (
            O => \N__31365\,
            I => \N__31362\
        );

    \I__5185\ : Span4Mux_h
    port map (
            O => \N__31362\,
            I => \N__31357\
        );

    \I__5184\ : InMux
    port map (
            O => \N__31361\,
            I => \N__31354\
        );

    \I__5183\ : InMux
    port map (
            O => \N__31360\,
            I => \N__31351\
        );

    \I__5182\ : Span4Mux_v
    port map (
            O => \N__31357\,
            I => \N__31345\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__31354\,
            I => \N__31345\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__31351\,
            I => \N__31342\
        );

    \I__5179\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31339\
        );

    \I__5178\ : Span4Mux_v
    port map (
            O => \N__31345\,
            I => \N__31336\
        );

    \I__5177\ : Odrv4
    port map (
            O => \N__31342\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__31339\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5175\ : Odrv4
    port map (
            O => \N__31336\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5174\ : InMux
    port map (
            O => \N__31329\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__5173\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31323\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__31323\,
            I => \N__31320\
        );

    \I__5171\ : Span4Mux_h
    port map (
            O => \N__31320\,
            I => \N__31317\
        );

    \I__5170\ : Span4Mux_h
    port map (
            O => \N__31317\,
            I => \N__31314\
        );

    \I__5169\ : Span4Mux_v
    port map (
            O => \N__31314\,
            I => \N__31311\
        );

    \I__5168\ : Odrv4
    port map (
            O => \N__31311\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__5167\ : CascadeMux
    port map (
            O => \N__31308\,
            I => \N__31304\
        );

    \I__5166\ : CascadeMux
    port map (
            O => \N__31307\,
            I => \N__31300\
        );

    \I__5165\ : InMux
    port map (
            O => \N__31304\,
            I => \N__31297\
        );

    \I__5164\ : InMux
    port map (
            O => \N__31303\,
            I => \N__31293\
        );

    \I__5163\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31290\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__31297\,
            I => \N__31287\
        );

    \I__5161\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31284\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__31293\,
            I => \N__31281\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__31290\,
            I => \N__31278\
        );

    \I__5158\ : Span12Mux_h
    port map (
            O => \N__31287\,
            I => \N__31275\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__31284\,
            I => \N__31272\
        );

    \I__5156\ : Span4Mux_v
    port map (
            O => \N__31281\,
            I => \N__31267\
        );

    \I__5155\ : Span4Mux_v
    port map (
            O => \N__31278\,
            I => \N__31267\
        );

    \I__5154\ : Odrv12
    port map (
            O => \N__31275\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__31272\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__5152\ : Odrv4
    port map (
            O => \N__31267\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__5151\ : InMux
    port map (
            O => \N__31260\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__5150\ : InMux
    port map (
            O => \N__31257\,
            I => \N__31254\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__31254\,
            I => \N__31251\
        );

    \I__5148\ : Span4Mux_h
    port map (
            O => \N__31251\,
            I => \N__31248\
        );

    \I__5147\ : Span4Mux_h
    port map (
            O => \N__31248\,
            I => \N__31245\
        );

    \I__5146\ : Odrv4
    port map (
            O => \N__31245\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__31242\,
            I => \N__31239\
        );

    \I__5144\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31236\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__31236\,
            I => \N__31233\
        );

    \I__5142\ : Span4Mux_v
    port map (
            O => \N__31233\,
            I => \N__31230\
        );

    \I__5141\ : Span4Mux_h
    port map (
            O => \N__31230\,
            I => \N__31224\
        );

    \I__5140\ : CascadeMux
    port map (
            O => \N__31229\,
            I => \N__31221\
        );

    \I__5139\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31218\
        );

    \I__5138\ : InMux
    port map (
            O => \N__31227\,
            I => \N__31215\
        );

    \I__5137\ : Span4Mux_h
    port map (
            O => \N__31224\,
            I => \N__31212\
        );

    \I__5136\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31209\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__31218\,
            I => \N__31206\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__31215\,
            I => \N__31203\
        );

    \I__5133\ : Span4Mux_v
    port map (
            O => \N__31212\,
            I => \N__31200\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__31209\,
            I => \N__31193\
        );

    \I__5131\ : Span4Mux_h
    port map (
            O => \N__31206\,
            I => \N__31193\
        );

    \I__5130\ : Span4Mux_h
    port map (
            O => \N__31203\,
            I => \N__31193\
        );

    \I__5129\ : Odrv4
    port map (
            O => \N__31200\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__31193\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__5127\ : InMux
    port map (
            O => \N__31188\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__5126\ : InMux
    port map (
            O => \N__31185\,
            I => \N__31182\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__31182\,
            I => \N__31179\
        );

    \I__5124\ : Span4Mux_v
    port map (
            O => \N__31179\,
            I => \N__31176\
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__31176\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__5122\ : CascadeMux
    port map (
            O => \N__31173\,
            I => \N__31170\
        );

    \I__5121\ : InMux
    port map (
            O => \N__31170\,
            I => \N__31167\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__31167\,
            I => \N__31164\
        );

    \I__5119\ : Span4Mux_h
    port map (
            O => \N__31164\,
            I => \N__31161\
        );

    \I__5118\ : Span4Mux_h
    port map (
            O => \N__31161\,
            I => \N__31158\
        );

    \I__5117\ : Span4Mux_v
    port map (
            O => \N__31158\,
            I => \N__31152\
        );

    \I__5116\ : InMux
    port map (
            O => \N__31157\,
            I => \N__31147\
        );

    \I__5115\ : InMux
    port map (
            O => \N__31156\,
            I => \N__31147\
        );

    \I__5114\ : InMux
    port map (
            O => \N__31155\,
            I => \N__31144\
        );

    \I__5113\ : Span4Mux_v
    port map (
            O => \N__31152\,
            I => \N__31139\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__31147\,
            I => \N__31139\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__31144\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__5110\ : Odrv4
    port map (
            O => \N__31139\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__5109\ : InMux
    port map (
            O => \N__31134\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__5108\ : InMux
    port map (
            O => \N__31131\,
            I => \N__31128\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__31128\,
            I => \N__31125\
        );

    \I__5106\ : Span12Mux_h
    port map (
            O => \N__31125\,
            I => \N__31122\
        );

    \I__5105\ : Odrv12
    port map (
            O => \N__31122\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__5104\ : CascadeMux
    port map (
            O => \N__31119\,
            I => \N__31116\
        );

    \I__5103\ : InMux
    port map (
            O => \N__31116\,
            I => \N__31111\
        );

    \I__5102\ : InMux
    port map (
            O => \N__31115\,
            I => \N__31108\
        );

    \I__5101\ : InMux
    port map (
            O => \N__31114\,
            I => \N__31105\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__31111\,
            I => \N__31102\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__31108\,
            I => \N__31098\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__31105\,
            I => \N__31095\
        );

    \I__5097\ : Span12Mux_v
    port map (
            O => \N__31102\,
            I => \N__31092\
        );

    \I__5096\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31089\
        );

    \I__5095\ : Span4Mux_h
    port map (
            O => \N__31098\,
            I => \N__31084\
        );

    \I__5094\ : Span4Mux_h
    port map (
            O => \N__31095\,
            I => \N__31084\
        );

    \I__5093\ : Odrv12
    port map (
            O => \N__31092\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__31089\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5091\ : Odrv4
    port map (
            O => \N__31084\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5090\ : InMux
    port map (
            O => \N__31077\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__5089\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31071\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__31071\,
            I => \N__31068\
        );

    \I__5087\ : Span4Mux_h
    port map (
            O => \N__31068\,
            I => \N__31065\
        );

    \I__5086\ : Odrv4
    port map (
            O => \N__31065\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__5085\ : CascadeMux
    port map (
            O => \N__31062\,
            I => \N__31059\
        );

    \I__5084\ : InMux
    port map (
            O => \N__31059\,
            I => \N__31056\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__31056\,
            I => \N__31053\
        );

    \I__5082\ : Span4Mux_v
    port map (
            O => \N__31053\,
            I => \N__31050\
        );

    \I__5081\ : Span4Mux_v
    port map (
            O => \N__31050\,
            I => \N__31046\
        );

    \I__5080\ : CascadeMux
    port map (
            O => \N__31049\,
            I => \N__31043\
        );

    \I__5079\ : Span4Mux_v
    port map (
            O => \N__31046\,
            I => \N__31038\
        );

    \I__5078\ : InMux
    port map (
            O => \N__31043\,
            I => \N__31033\
        );

    \I__5077\ : InMux
    port map (
            O => \N__31042\,
            I => \N__31033\
        );

    \I__5076\ : InMux
    port map (
            O => \N__31041\,
            I => \N__31030\
        );

    \I__5075\ : Span4Mux_h
    port map (
            O => \N__31038\,
            I => \N__31025\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__31033\,
            I => \N__31025\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__31030\,
            I => \N__31020\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__31025\,
            I => \N__31020\
        );

    \I__5071\ : Odrv4
    port map (
            O => \N__31020\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5070\ : InMux
    port map (
            O => \N__31017\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__5069\ : InMux
    port map (
            O => \N__31014\,
            I => \N__31011\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__31011\,
            I => \N__31008\
        );

    \I__5067\ : Span4Mux_h
    port map (
            O => \N__31008\,
            I => \N__31005\
        );

    \I__5066\ : Span4Mux_h
    port map (
            O => \N__31005\,
            I => \N__31002\
        );

    \I__5065\ : Odrv4
    port map (
            O => \N__31002\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__5064\ : CascadeMux
    port map (
            O => \N__30999\,
            I => \N__30996\
        );

    \I__5063\ : InMux
    port map (
            O => \N__30996\,
            I => \N__30993\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__30993\,
            I => \N__30990\
        );

    \I__5061\ : Span4Mux_v
    port map (
            O => \N__30990\,
            I => \N__30986\
        );

    \I__5060\ : CascadeMux
    port map (
            O => \N__30989\,
            I => \N__30983\
        );

    \I__5059\ : Sp12to4
    port map (
            O => \N__30986\,
            I => \N__30978\
        );

    \I__5058\ : InMux
    port map (
            O => \N__30983\,
            I => \N__30973\
        );

    \I__5057\ : InMux
    port map (
            O => \N__30982\,
            I => \N__30973\
        );

    \I__5056\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30970\
        );

    \I__5055\ : Span12Mux_h
    port map (
            O => \N__30978\,
            I => \N__30967\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__30973\,
            I => \N__30964\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__30970\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__5052\ : Odrv12
    port map (
            O => \N__30967\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__30964\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__5050\ : InMux
    port map (
            O => \N__30957\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\
        );

    \I__5049\ : InMux
    port map (
            O => \N__30954\,
            I => \N__30951\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__30951\,
            I => \N__30948\
        );

    \I__5047\ : Span4Mux_h
    port map (
            O => \N__30948\,
            I => \N__30945\
        );

    \I__5046\ : Odrv4
    port map (
            O => \N__30945\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__5045\ : CascadeMux
    port map (
            O => \N__30942\,
            I => \N__30939\
        );

    \I__5044\ : InMux
    port map (
            O => \N__30939\,
            I => \N__30936\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__30936\,
            I => \N__30933\
        );

    \I__5042\ : Span4Mux_h
    port map (
            O => \N__30933\,
            I => \N__30930\
        );

    \I__5041\ : Span4Mux_h
    port map (
            O => \N__30930\,
            I => \N__30924\
        );

    \I__5040\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30921\
        );

    \I__5039\ : CascadeMux
    port map (
            O => \N__30928\,
            I => \N__30918\
        );

    \I__5038\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30915\
        );

    \I__5037\ : Sp12to4
    port map (
            O => \N__30924\,
            I => \N__30910\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__30921\,
            I => \N__30910\
        );

    \I__5035\ : InMux
    port map (
            O => \N__30918\,
            I => \N__30907\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__30915\,
            I => \N__30904\
        );

    \I__5033\ : Span12Mux_v
    port map (
            O => \N__30910\,
            I => \N__30901\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__30907\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__5031\ : Odrv4
    port map (
            O => \N__30904\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__5030\ : Odrv12
    port map (
            O => \N__30901\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__5029\ : InMux
    port map (
            O => \N__30894\,
            I => \bfn_11_20_0_\
        );

    \I__5028\ : InMux
    port map (
            O => \N__30891\,
            I => \N__30888\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__30888\,
            I => \N__30885\
        );

    \I__5026\ : Span4Mux_h
    port map (
            O => \N__30885\,
            I => \N__30882\
        );

    \I__5025\ : Span4Mux_h
    port map (
            O => \N__30882\,
            I => \N__30879\
        );

    \I__5024\ : Span4Mux_v
    port map (
            O => \N__30879\,
            I => \N__30876\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__30876\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__5022\ : CascadeMux
    port map (
            O => \N__30873\,
            I => \N__30870\
        );

    \I__5021\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30867\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__30867\,
            I => \N__30864\
        );

    \I__5019\ : Span4Mux_v
    port map (
            O => \N__30864\,
            I => \N__30861\
        );

    \I__5018\ : Span4Mux_h
    port map (
            O => \N__30861\,
            I => \N__30857\
        );

    \I__5017\ : CascadeMux
    port map (
            O => \N__30860\,
            I => \N__30854\
        );

    \I__5016\ : Span4Mux_h
    port map (
            O => \N__30857\,
            I => \N__30849\
        );

    \I__5015\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30846\
        );

    \I__5014\ : InMux
    port map (
            O => \N__30853\,
            I => \N__30843\
        );

    \I__5013\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30840\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__30849\,
            I => \N__30835\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__30846\,
            I => \N__30835\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__30843\,
            I => \N__30830\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__30840\,
            I => \N__30830\
        );

    \I__5008\ : Odrv4
    port map (
            O => \N__30835\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__30830\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__5006\ : InMux
    port map (
            O => \N__30825\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__5005\ : InMux
    port map (
            O => \N__30822\,
            I => \N__30819\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__30819\,
            I => \N__30816\
        );

    \I__5003\ : Span4Mux_v
    port map (
            O => \N__30816\,
            I => \N__30813\
        );

    \I__5002\ : Span4Mux_v
    port map (
            O => \N__30813\,
            I => \N__30810\
        );

    \I__5001\ : Odrv4
    port map (
            O => \N__30810\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__5000\ : CascadeMux
    port map (
            O => \N__30807\,
            I => \N__30804\
        );

    \I__4999\ : InMux
    port map (
            O => \N__30804\,
            I => \N__30801\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__30801\,
            I => \N__30798\
        );

    \I__4997\ : Span4Mux_h
    port map (
            O => \N__30798\,
            I => \N__30795\
        );

    \I__4996\ : Span4Mux_h
    port map (
            O => \N__30795\,
            I => \N__30790\
        );

    \I__4995\ : CascadeMux
    port map (
            O => \N__30794\,
            I => \N__30787\
        );

    \I__4994\ : InMux
    port map (
            O => \N__30793\,
            I => \N__30784\
        );

    \I__4993\ : Span4Mux_v
    port map (
            O => \N__30790\,
            I => \N__30781\
        );

    \I__4992\ : InMux
    port map (
            O => \N__30787\,
            I => \N__30778\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__30784\,
            I => \N__30775\
        );

    \I__4990\ : Span4Mux_v
    port map (
            O => \N__30781\,
            I => \N__30771\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__30778\,
            I => \N__30766\
        );

    \I__4988\ : Span4Mux_h
    port map (
            O => \N__30775\,
            I => \N__30766\
        );

    \I__4987\ : InMux
    port map (
            O => \N__30774\,
            I => \N__30763\
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__30771\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__4985\ : Odrv4
    port map (
            O => \N__30766\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__30763\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__4983\ : InMux
    port map (
            O => \N__30756\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__4982\ : InMux
    port map (
            O => \N__30753\,
            I => \N__30750\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__30750\,
            I => \N__30747\
        );

    \I__4980\ : Span4Mux_v
    port map (
            O => \N__30747\,
            I => \N__30744\
        );

    \I__4979\ : Span4Mux_h
    port map (
            O => \N__30744\,
            I => \N__30741\
        );

    \I__4978\ : Odrv4
    port map (
            O => \N__30741\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__4977\ : CascadeMux
    port map (
            O => \N__30738\,
            I => \N__30735\
        );

    \I__4976\ : InMux
    port map (
            O => \N__30735\,
            I => \N__30732\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__30732\,
            I => \N__30728\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__30731\,
            I => \N__30724\
        );

    \I__4973\ : Span4Mux_v
    port map (
            O => \N__30728\,
            I => \N__30720\
        );

    \I__4972\ : InMux
    port map (
            O => \N__30727\,
            I => \N__30717\
        );

    \I__4971\ : InMux
    port map (
            O => \N__30724\,
            I => \N__30714\
        );

    \I__4970\ : InMux
    port map (
            O => \N__30723\,
            I => \N__30711\
        );

    \I__4969\ : Span4Mux_h
    port map (
            O => \N__30720\,
            I => \N__30708\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__30717\,
            I => \N__30705\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__30714\,
            I => \N__30702\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__30711\,
            I => \N__30699\
        );

    \I__4965\ : Span4Mux_h
    port map (
            O => \N__30708\,
            I => \N__30694\
        );

    \I__4964\ : Span4Mux_h
    port map (
            O => \N__30705\,
            I => \N__30694\
        );

    \I__4963\ : Odrv12
    port map (
            O => \N__30702\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4962\ : Odrv4
    port map (
            O => \N__30699\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4961\ : Odrv4
    port map (
            O => \N__30694\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4960\ : InMux
    port map (
            O => \N__30687\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__4959\ : InMux
    port map (
            O => \N__30684\,
            I => \N__30681\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__30681\,
            I => \N__30678\
        );

    \I__4957\ : Span4Mux_v
    port map (
            O => \N__30678\,
            I => \N__30675\
        );

    \I__4956\ : Span4Mux_v
    port map (
            O => \N__30675\,
            I => \N__30672\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__30672\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__4954\ : CascadeMux
    port map (
            O => \N__30669\,
            I => \N__30666\
        );

    \I__4953\ : InMux
    port map (
            O => \N__30666\,
            I => \N__30663\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__30663\,
            I => \N__30660\
        );

    \I__4951\ : Span4Mux_v
    port map (
            O => \N__30660\,
            I => \N__30657\
        );

    \I__4950\ : Sp12to4
    port map (
            O => \N__30657\,
            I => \N__30652\
        );

    \I__4949\ : InMux
    port map (
            O => \N__30656\,
            I => \N__30648\
        );

    \I__4948\ : InMux
    port map (
            O => \N__30655\,
            I => \N__30645\
        );

    \I__4947\ : Span12Mux_h
    port map (
            O => \N__30652\,
            I => \N__30642\
        );

    \I__4946\ : InMux
    port map (
            O => \N__30651\,
            I => \N__30639\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__30648\,
            I => \N__30636\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__30645\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__4943\ : Odrv12
    port map (
            O => \N__30642\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__30639\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__4941\ : Odrv4
    port map (
            O => \N__30636\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__4940\ : InMux
    port map (
            O => \N__30627\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__4939\ : InMux
    port map (
            O => \N__30624\,
            I => \N__30621\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__30621\,
            I => \N__30618\
        );

    \I__4937\ : Span4Mux_v
    port map (
            O => \N__30618\,
            I => \N__30615\
        );

    \I__4936\ : Span4Mux_h
    port map (
            O => \N__30615\,
            I => \N__30612\
        );

    \I__4935\ : Odrv4
    port map (
            O => \N__30612\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__4934\ : CascadeMux
    port map (
            O => \N__30609\,
            I => \N__30606\
        );

    \I__4933\ : InMux
    port map (
            O => \N__30606\,
            I => \N__30603\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__30603\,
            I => \N__30599\
        );

    \I__4931\ : InMux
    port map (
            O => \N__30602\,
            I => \N__30594\
        );

    \I__4930\ : Span12Mux_v
    port map (
            O => \N__30599\,
            I => \N__30591\
        );

    \I__4929\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30588\
        );

    \I__4928\ : InMux
    port map (
            O => \N__30597\,
            I => \N__30585\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__30594\,
            I => \N__30582\
        );

    \I__4926\ : Odrv12
    port map (
            O => \N__30591\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__30588\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__30585\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__30582\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4922\ : InMux
    port map (
            O => \N__30573\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__4921\ : InMux
    port map (
            O => \N__30570\,
            I => \N__30567\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__30567\,
            I => \N__30564\
        );

    \I__4919\ : Span4Mux_v
    port map (
            O => \N__30564\,
            I => \N__30561\
        );

    \I__4918\ : Span4Mux_v
    port map (
            O => \N__30561\,
            I => \N__30558\
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__30558\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__4916\ : CascadeMux
    port map (
            O => \N__30555\,
            I => \N__30552\
        );

    \I__4915\ : InMux
    port map (
            O => \N__30552\,
            I => \N__30549\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__30549\,
            I => \N__30544\
        );

    \I__4913\ : CascadeMux
    port map (
            O => \N__30548\,
            I => \N__30541\
        );

    \I__4912\ : InMux
    port map (
            O => \N__30547\,
            I => \N__30537\
        );

    \I__4911\ : Span4Mux_v
    port map (
            O => \N__30544\,
            I => \N__30534\
        );

    \I__4910\ : InMux
    port map (
            O => \N__30541\,
            I => \N__30531\
        );

    \I__4909\ : InMux
    port map (
            O => \N__30540\,
            I => \N__30528\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__30537\,
            I => \N__30525\
        );

    \I__4907\ : Span4Mux_h
    port map (
            O => \N__30534\,
            I => \N__30522\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__30531\,
            I => \N__30519\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__30528\,
            I => \N__30516\
        );

    \I__4904\ : Span4Mux_v
    port map (
            O => \N__30525\,
            I => \N__30513\
        );

    \I__4903\ : Span4Mux_h
    port map (
            O => \N__30522\,
            I => \N__30508\
        );

    \I__4902\ : Span4Mux_v
    port map (
            O => \N__30519\,
            I => \N__30508\
        );

    \I__4901\ : Span4Mux_v
    port map (
            O => \N__30516\,
            I => \N__30505\
        );

    \I__4900\ : Odrv4
    port map (
            O => \N__30513\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4899\ : Odrv4
    port map (
            O => \N__30508\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4898\ : Odrv4
    port map (
            O => \N__30505\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4897\ : InMux
    port map (
            O => \N__30498\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__4896\ : InMux
    port map (
            O => \N__30495\,
            I => \N__30492\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__30492\,
            I => \N__30489\
        );

    \I__4894\ : Span12Mux_v
    port map (
            O => \N__30489\,
            I => \N__30486\
        );

    \I__4893\ : Odrv12
    port map (
            O => \N__30486\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__4892\ : CascadeMux
    port map (
            O => \N__30483\,
            I => \N__30479\
        );

    \I__4891\ : CascadeMux
    port map (
            O => \N__30482\,
            I => \N__30475\
        );

    \I__4890\ : InMux
    port map (
            O => \N__30479\,
            I => \N__30472\
        );

    \I__4889\ : InMux
    port map (
            O => \N__30478\,
            I => \N__30469\
        );

    \I__4888\ : InMux
    port map (
            O => \N__30475\,
            I => \N__30466\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__30472\,
            I => \N__30463\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__30469\,
            I => \N__30459\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__30466\,
            I => \N__30456\
        );

    \I__4884\ : Span12Mux_v
    port map (
            O => \N__30463\,
            I => \N__30453\
        );

    \I__4883\ : InMux
    port map (
            O => \N__30462\,
            I => \N__30450\
        );

    \I__4882\ : Span4Mux_v
    port map (
            O => \N__30459\,
            I => \N__30445\
        );

    \I__4881\ : Span4Mux_h
    port map (
            O => \N__30456\,
            I => \N__30445\
        );

    \I__4880\ : Odrv12
    port map (
            O => \N__30453\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__30450\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__4878\ : Odrv4
    port map (
            O => \N__30445\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__4877\ : InMux
    port map (
            O => \N__30438\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\
        );

    \I__4876\ : InMux
    port map (
            O => \N__30435\,
            I => \N__30432\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__30432\,
            I => \N__30428\
        );

    \I__4874\ : InMux
    port map (
            O => \N__30431\,
            I => \N__30424\
        );

    \I__4873\ : Span12Mux_h
    port map (
            O => \N__30428\,
            I => \N__30421\
        );

    \I__4872\ : InMux
    port map (
            O => \N__30427\,
            I => \N__30418\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__30424\,
            I => \N__30415\
        );

    \I__4870\ : Odrv12
    port map (
            O => \N__30421\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__30418\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4868\ : Odrv4
    port map (
            O => \N__30415\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4867\ : CascadeMux
    port map (
            O => \N__30408\,
            I => \N__30405\
        );

    \I__4866\ : InMux
    port map (
            O => \N__30405\,
            I => \N__30402\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__30402\,
            I => \N__30399\
        );

    \I__4864\ : Span4Mux_h
    port map (
            O => \N__30399\,
            I => \N__30396\
        );

    \I__4863\ : Odrv4
    port map (
            O => \N__30396\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__4862\ : InMux
    port map (
            O => \N__30393\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__4861\ : InMux
    port map (
            O => \N__30390\,
            I => \N__30387\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__30387\,
            I => \N__30384\
        );

    \I__4859\ : Span4Mux_h
    port map (
            O => \N__30384\,
            I => \N__30381\
        );

    \I__4858\ : Span4Mux_h
    port map (
            O => \N__30381\,
            I => \N__30378\
        );

    \I__4857\ : Odrv4
    port map (
            O => \N__30378\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__4856\ : CascadeMux
    port map (
            O => \N__30375\,
            I => \N__30372\
        );

    \I__4855\ : InMux
    port map (
            O => \N__30372\,
            I => \N__30369\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__30369\,
            I => \N__30365\
        );

    \I__4853\ : CascadeMux
    port map (
            O => \N__30368\,
            I => \N__30362\
        );

    \I__4852\ : Span4Mux_v
    port map (
            O => \N__30365\,
            I => \N__30359\
        );

    \I__4851\ : InMux
    port map (
            O => \N__30362\,
            I => \N__30356\
        );

    \I__4850\ : Span4Mux_h
    port map (
            O => \N__30359\,
            I => \N__30353\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__30356\,
            I => \N__30348\
        );

    \I__4848\ : Span4Mux_h
    port map (
            O => \N__30353\,
            I => \N__30345\
        );

    \I__4847\ : InMux
    port map (
            O => \N__30352\,
            I => \N__30342\
        );

    \I__4846\ : InMux
    port map (
            O => \N__30351\,
            I => \N__30339\
        );

    \I__4845\ : Span4Mux_h
    port map (
            O => \N__30348\,
            I => \N__30334\
        );

    \I__4844\ : Span4Mux_v
    port map (
            O => \N__30345\,
            I => \N__30334\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__30342\,
            I => \N__30331\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__30339\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__30334\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__4840\ : Odrv4
    port map (
            O => \N__30331\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__4839\ : InMux
    port map (
            O => \N__30324\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__4838\ : InMux
    port map (
            O => \N__30321\,
            I => \N__30318\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__30318\,
            I => \N__30315\
        );

    \I__4836\ : Span4Mux_v
    port map (
            O => \N__30315\,
            I => \N__30312\
        );

    \I__4835\ : Odrv4
    port map (
            O => \N__30312\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__4834\ : CascadeMux
    port map (
            O => \N__30309\,
            I => \N__30306\
        );

    \I__4833\ : InMux
    port map (
            O => \N__30306\,
            I => \N__30303\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__30303\,
            I => \N__30300\
        );

    \I__4831\ : Span4Mux_v
    port map (
            O => \N__30300\,
            I => \N__30297\
        );

    \I__4830\ : Sp12to4
    port map (
            O => \N__30297\,
            I => \N__30291\
        );

    \I__4829\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30288\
        );

    \I__4828\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30285\
        );

    \I__4827\ : InMux
    port map (
            O => \N__30294\,
            I => \N__30282\
        );

    \I__4826\ : Span12Mux_h
    port map (
            O => \N__30291\,
            I => \N__30279\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__30288\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__30285\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__30282\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__4822\ : Odrv12
    port map (
            O => \N__30279\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__4821\ : InMux
    port map (
            O => \N__30270\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__4820\ : InMux
    port map (
            O => \N__30267\,
            I => \N__30264\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__30264\,
            I => \N__30261\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__30261\,
            I => \N__30258\
        );

    \I__4817\ : Span4Mux_v
    port map (
            O => \N__30258\,
            I => \N__30255\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__30255\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__4815\ : CascadeMux
    port map (
            O => \N__30252\,
            I => \N__30249\
        );

    \I__4814\ : InMux
    port map (
            O => \N__30249\,
            I => \N__30246\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__30246\,
            I => \N__30243\
        );

    \I__4812\ : Span4Mux_h
    port map (
            O => \N__30243\,
            I => \N__30240\
        );

    \I__4811\ : Span4Mux_h
    port map (
            O => \N__30240\,
            I => \N__30236\
        );

    \I__4810\ : InMux
    port map (
            O => \N__30239\,
            I => \N__30233\
        );

    \I__4809\ : Span4Mux_h
    port map (
            O => \N__30236\,
            I => \N__30229\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__30233\,
            I => \N__30225\
        );

    \I__4807\ : InMux
    port map (
            O => \N__30232\,
            I => \N__30222\
        );

    \I__4806\ : Sp12to4
    port map (
            O => \N__30229\,
            I => \N__30219\
        );

    \I__4805\ : InMux
    port map (
            O => \N__30228\,
            I => \N__30216\
        );

    \I__4804\ : Span4Mux_h
    port map (
            O => \N__30225\,
            I => \N__30213\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__30222\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__4802\ : Odrv12
    port map (
            O => \N__30219\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__30216\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__4800\ : Odrv4
    port map (
            O => \N__30213\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__4799\ : InMux
    port map (
            O => \N__30204\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__4798\ : InMux
    port map (
            O => \N__30201\,
            I => \N__30198\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__30198\,
            I => \N__30195\
        );

    \I__4796\ : Span4Mux_v
    port map (
            O => \N__30195\,
            I => \N__30192\
        );

    \I__4795\ : Span4Mux_v
    port map (
            O => \N__30192\,
            I => \N__30189\
        );

    \I__4794\ : Odrv4
    port map (
            O => \N__30189\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__4793\ : CascadeMux
    port map (
            O => \N__30186\,
            I => \N__30183\
        );

    \I__4792\ : InMux
    port map (
            O => \N__30183\,
            I => \N__30180\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__30180\,
            I => \N__30177\
        );

    \I__4790\ : Span4Mux_v
    port map (
            O => \N__30177\,
            I => \N__30174\
        );

    \I__4789\ : Sp12to4
    port map (
            O => \N__30174\,
            I => \N__30168\
        );

    \I__4788\ : InMux
    port map (
            O => \N__30173\,
            I => \N__30165\
        );

    \I__4787\ : InMux
    port map (
            O => \N__30172\,
            I => \N__30162\
        );

    \I__4786\ : InMux
    port map (
            O => \N__30171\,
            I => \N__30159\
        );

    \I__4785\ : Span12Mux_h
    port map (
            O => \N__30168\,
            I => \N__30156\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__30165\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__30162\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__30159\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4781\ : Odrv12
    port map (
            O => \N__30156\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4780\ : InMux
    port map (
            O => \N__30147\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__4779\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30141\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__30141\,
            I => \N__30138\
        );

    \I__4777\ : Span4Mux_v
    port map (
            O => \N__30138\,
            I => \N__30135\
        );

    \I__4776\ : Span4Mux_h
    port map (
            O => \N__30135\,
            I => \N__30132\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__30132\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__4774\ : CascadeMux
    port map (
            O => \N__30129\,
            I => \N__30126\
        );

    \I__4773\ : InMux
    port map (
            O => \N__30126\,
            I => \N__30123\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__30123\,
            I => \N__30120\
        );

    \I__4771\ : Span4Mux_v
    port map (
            O => \N__30120\,
            I => \N__30117\
        );

    \I__4770\ : Span4Mux_h
    port map (
            O => \N__30117\,
            I => \N__30114\
        );

    \I__4769\ : Span4Mux_h
    port map (
            O => \N__30114\,
            I => \N__30110\
        );

    \I__4768\ : InMux
    port map (
            O => \N__30113\,
            I => \N__30107\
        );

    \I__4767\ : Span4Mux_v
    port map (
            O => \N__30110\,
            I => \N__30100\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__30107\,
            I => \N__30100\
        );

    \I__4765\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30097\
        );

    \I__4764\ : InMux
    port map (
            O => \N__30105\,
            I => \N__30094\
        );

    \I__4763\ : Span4Mux_v
    port map (
            O => \N__30100\,
            I => \N__30091\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__30097\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__30094\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__4760\ : Odrv4
    port map (
            O => \N__30091\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__4759\ : InMux
    port map (
            O => \N__30084\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__4758\ : InMux
    port map (
            O => \N__30081\,
            I => \N__30078\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__30078\,
            I => \N__30075\
        );

    \I__4756\ : Odrv12
    port map (
            O => \N__30075\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__4755\ : CascadeMux
    port map (
            O => \N__30072\,
            I => \N__30069\
        );

    \I__4754\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30066\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__30066\,
            I => \N__30063\
        );

    \I__4752\ : Span4Mux_v
    port map (
            O => \N__30063\,
            I => \N__30060\
        );

    \I__4751\ : Sp12to4
    port map (
            O => \N__30060\,
            I => \N__30054\
        );

    \I__4750\ : InMux
    port map (
            O => \N__30059\,
            I => \N__30051\
        );

    \I__4749\ : InMux
    port map (
            O => \N__30058\,
            I => \N__30048\
        );

    \I__4748\ : InMux
    port map (
            O => \N__30057\,
            I => \N__30045\
        );

    \I__4747\ : Span12Mux_v
    port map (
            O => \N__30054\,
            I => \N__30042\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__30051\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__30048\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__30045\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__4743\ : Odrv12
    port map (
            O => \N__30042\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__4742\ : InMux
    port map (
            O => \N__30033\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\
        );

    \I__4741\ : CascadeMux
    port map (
            O => \N__30030\,
            I => \N__30027\
        );

    \I__4740\ : InMux
    port map (
            O => \N__30027\,
            I => \N__30024\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__30024\,
            I => \N__30019\
        );

    \I__4738\ : InMux
    port map (
            O => \N__30023\,
            I => \N__30016\
        );

    \I__4737\ : InMux
    port map (
            O => \N__30022\,
            I => \N__30013\
        );

    \I__4736\ : Span4Mux_v
    port map (
            O => \N__30019\,
            I => \N__30008\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__30016\,
            I => \N__30008\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__30013\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__4733\ : Odrv4
    port map (
            O => \N__30008\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__4732\ : InMux
    port map (
            O => \N__30003\,
            I => \bfn_11_18_0_\
        );

    \I__4731\ : InMux
    port map (
            O => \N__30000\,
            I => \N__29997\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__29997\,
            I => \N__29994\
        );

    \I__4729\ : Span4Mux_h
    port map (
            O => \N__29994\,
            I => \N__29991\
        );

    \I__4728\ : Span4Mux_v
    port map (
            O => \N__29991\,
            I => \N__29988\
        );

    \I__4727\ : Odrv4
    port map (
            O => \N__29988\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__4726\ : InMux
    port map (
            O => \N__29985\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__4725\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29979\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__29979\,
            I => \N__29975\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__29978\,
            I => \N__29972\
        );

    \I__4722\ : Span4Mux_h
    port map (
            O => \N__29975\,
            I => \N__29968\
        );

    \I__4721\ : InMux
    port map (
            O => \N__29972\,
            I => \N__29965\
        );

    \I__4720\ : InMux
    port map (
            O => \N__29971\,
            I => \N__29962\
        );

    \I__4719\ : Odrv4
    port map (
            O => \N__29968\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__29965\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__29962\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__4716\ : InMux
    port map (
            O => \N__29955\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__4715\ : InMux
    port map (
            O => \N__29952\,
            I => \N__29949\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__29949\,
            I => \N__29946\
        );

    \I__4713\ : Span4Mux_h
    port map (
            O => \N__29946\,
            I => \N__29941\
        );

    \I__4712\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29938\
        );

    \I__4711\ : InMux
    port map (
            O => \N__29944\,
            I => \N__29935\
        );

    \I__4710\ : Span4Mux_v
    port map (
            O => \N__29941\,
            I => \N__29930\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__29938\,
            I => \N__29930\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__29935\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__4707\ : Odrv4
    port map (
            O => \N__29930\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__4706\ : InMux
    port map (
            O => \N__29925\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__4705\ : InMux
    port map (
            O => \N__29922\,
            I => \N__29918\
        );

    \I__4704\ : InMux
    port map (
            O => \N__29921\,
            I => \N__29914\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__29918\,
            I => \N__29911\
        );

    \I__4702\ : InMux
    port map (
            O => \N__29917\,
            I => \N__29908\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__29914\,
            I => \N__29905\
        );

    \I__4700\ : Span4Mux_v
    port map (
            O => \N__29911\,
            I => \N__29900\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__29908\,
            I => \N__29900\
        );

    \I__4698\ : Odrv12
    port map (
            O => \N__29905\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__4697\ : Odrv4
    port map (
            O => \N__29900\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__4696\ : InMux
    port map (
            O => \N__29895\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__4695\ : InMux
    port map (
            O => \N__29892\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__29889\,
            I => \N__29885\
        );

    \I__4693\ : InMux
    port map (
            O => \N__29888\,
            I => \N__29882\
        );

    \I__4692\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29876\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__29882\,
            I => \N__29873\
        );

    \I__4690\ : CascadeMux
    port map (
            O => \N__29881\,
            I => \N__29870\
        );

    \I__4689\ : InMux
    port map (
            O => \N__29880\,
            I => \N__29865\
        );

    \I__4688\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29865\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__29876\,
            I => \N__29860\
        );

    \I__4686\ : Span4Mux_v
    port map (
            O => \N__29873\,
            I => \N__29860\
        );

    \I__4685\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29857\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__29865\,
            I => \N__29854\
        );

    \I__4683\ : Sp12to4
    port map (
            O => \N__29860\,
            I => \N__29849\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__29857\,
            I => \N__29849\
        );

    \I__4681\ : Span12Mux_v
    port map (
            O => \N__29854\,
            I => \N__29844\
        );

    \I__4680\ : Span12Mux_h
    port map (
            O => \N__29849\,
            I => \N__29844\
        );

    \I__4679\ : Odrv12
    port map (
            O => \N__29844\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__4678\ : CascadeMux
    port map (
            O => \N__29841\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\
        );

    \I__4677\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29835\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__29835\,
            I => \N__29832\
        );

    \I__4675\ : Span4Mux_v
    port map (
            O => \N__29832\,
            I => \N__29829\
        );

    \I__4674\ : Odrv4
    port map (
            O => \N__29829\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__4673\ : InMux
    port map (
            O => \N__29826\,
            I => \N__29823\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__29823\,
            I => \N__29819\
        );

    \I__4671\ : InMux
    port map (
            O => \N__29822\,
            I => \N__29815\
        );

    \I__4670\ : Span4Mux_h
    port map (
            O => \N__29819\,
            I => \N__29812\
        );

    \I__4669\ : InMux
    port map (
            O => \N__29818\,
            I => \N__29809\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__29815\,
            I => \N__29806\
        );

    \I__4667\ : Odrv4
    port map (
            O => \N__29812\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__29809\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__4665\ : Odrv4
    port map (
            O => \N__29806\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__29799\,
            I => \N__29796\
        );

    \I__4663\ : InMux
    port map (
            O => \N__29796\,
            I => \N__29793\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__29793\,
            I => \N__29790\
        );

    \I__4661\ : Span4Mux_h
    port map (
            O => \N__29790\,
            I => \N__29787\
        );

    \I__4660\ : Odrv4
    port map (
            O => \N__29787\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__4659\ : InMux
    port map (
            O => \N__29784\,
            I => \N__29781\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__29781\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__4657\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29775\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__29775\,
            I => \N__29771\
        );

    \I__4655\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29767\
        );

    \I__4654\ : Span4Mux_h
    port map (
            O => \N__29771\,
            I => \N__29764\
        );

    \I__4653\ : InMux
    port map (
            O => \N__29770\,
            I => \N__29761\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__29767\,
            I => \N__29758\
        );

    \I__4651\ : Odrv4
    port map (
            O => \N__29764\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__29761\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__4649\ : Odrv4
    port map (
            O => \N__29758\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__4648\ : InMux
    port map (
            O => \N__29751\,
            I => \bfn_11_17_0_\
        );

    \I__4647\ : InMux
    port map (
            O => \N__29748\,
            I => \N__29745\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__29745\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__4645\ : InMux
    port map (
            O => \N__29742\,
            I => \N__29739\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__29739\,
            I => \N__29735\
        );

    \I__4643\ : InMux
    port map (
            O => \N__29738\,
            I => \N__29732\
        );

    \I__4642\ : Span4Mux_v
    port map (
            O => \N__29735\,
            I => \N__29728\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__29732\,
            I => \N__29725\
        );

    \I__4640\ : InMux
    port map (
            O => \N__29731\,
            I => \N__29722\
        );

    \I__4639\ : Span4Mux_h
    port map (
            O => \N__29728\,
            I => \N__29717\
        );

    \I__4638\ : Span4Mux_h
    port map (
            O => \N__29725\,
            I => \N__29717\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__29722\,
            I => \N__29714\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__29717\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__4635\ : Odrv4
    port map (
            O => \N__29714\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__4634\ : InMux
    port map (
            O => \N__29709\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__4633\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29703\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__29703\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__4631\ : InMux
    port map (
            O => \N__29700\,
            I => \N__29696\
        );

    \I__4630\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29693\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__29696\,
            I => \N__29690\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__29693\,
            I => \N__29686\
        );

    \I__4627\ : Span4Mux_h
    port map (
            O => \N__29690\,
            I => \N__29683\
        );

    \I__4626\ : InMux
    port map (
            O => \N__29689\,
            I => \N__29680\
        );

    \I__4625\ : Span4Mux_h
    port map (
            O => \N__29686\,
            I => \N__29677\
        );

    \I__4624\ : Span4Mux_v
    port map (
            O => \N__29683\,
            I => \N__29672\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__29680\,
            I => \N__29672\
        );

    \I__4622\ : Odrv4
    port map (
            O => \N__29677\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__4621\ : Odrv4
    port map (
            O => \N__29672\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__4620\ : InMux
    port map (
            O => \N__29667\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__4619\ : InMux
    port map (
            O => \N__29664\,
            I => \N__29661\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__29661\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__4617\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29654\
        );

    \I__4616\ : CascadeMux
    port map (
            O => \N__29657\,
            I => \N__29651\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__29654\,
            I => \N__29647\
        );

    \I__4614\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29644\
        );

    \I__4613\ : InMux
    port map (
            O => \N__29650\,
            I => \N__29641\
        );

    \I__4612\ : Span4Mux_h
    port map (
            O => \N__29647\,
            I => \N__29636\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__29644\,
            I => \N__29636\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__29641\,
            I => \N__29633\
        );

    \I__4609\ : Odrv4
    port map (
            O => \N__29636\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__4608\ : Odrv4
    port map (
            O => \N__29633\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__4607\ : InMux
    port map (
            O => \N__29628\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__4606\ : InMux
    port map (
            O => \N__29625\,
            I => \N__29622\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__29622\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__4604\ : CascadeMux
    port map (
            O => \N__29619\,
            I => \N__29615\
        );

    \I__4603\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29612\
        );

    \I__4602\ : InMux
    port map (
            O => \N__29615\,
            I => \N__29608\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__29612\,
            I => \N__29605\
        );

    \I__4600\ : InMux
    port map (
            O => \N__29611\,
            I => \N__29602\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__29608\,
            I => \N__29599\
        );

    \I__4598\ : Span4Mux_v
    port map (
            O => \N__29605\,
            I => \N__29594\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__29602\,
            I => \N__29594\
        );

    \I__4596\ : Odrv4
    port map (
            O => \N__29599\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__29594\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__4594\ : InMux
    port map (
            O => \N__29589\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__4593\ : InMux
    port map (
            O => \N__29586\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__4592\ : InMux
    port map (
            O => \N__29583\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__29580\,
            I => \N__29577\
        );

    \I__4590\ : InMux
    port map (
            O => \N__29577\,
            I => \N__29573\
        );

    \I__4589\ : InMux
    port map (
            O => \N__29576\,
            I => \N__29570\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__29573\,
            I => \N__29567\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__29570\,
            I => \N__29563\
        );

    \I__4586\ : Span4Mux_v
    port map (
            O => \N__29567\,
            I => \N__29560\
        );

    \I__4585\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29557\
        );

    \I__4584\ : Odrv12
    port map (
            O => \N__29563\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__29560\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__29557\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__4581\ : InMux
    port map (
            O => \N__29550\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__4580\ : CascadeMux
    port map (
            O => \N__29547\,
            I => \N__29544\
        );

    \I__4579\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29541\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__29541\,
            I => \N__29538\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__29538\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__4576\ : InMux
    port map (
            O => \N__29535\,
            I => \N__29531\
        );

    \I__4575\ : InMux
    port map (
            O => \N__29534\,
            I => \N__29528\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__29531\,
            I => \N__29524\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__29528\,
            I => \N__29521\
        );

    \I__4572\ : InMux
    port map (
            O => \N__29527\,
            I => \N__29518\
        );

    \I__4571\ : Span4Mux_v
    port map (
            O => \N__29524\,
            I => \N__29511\
        );

    \I__4570\ : Span4Mux_v
    port map (
            O => \N__29521\,
            I => \N__29511\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__29518\,
            I => \N__29511\
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__29511\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__4567\ : InMux
    port map (
            O => \N__29508\,
            I => \bfn_11_16_0_\
        );

    \I__4566\ : InMux
    port map (
            O => \N__29505\,
            I => \N__29502\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__29502\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__4564\ : InMux
    port map (
            O => \N__29499\,
            I => \N__29495\
        );

    \I__4563\ : InMux
    port map (
            O => \N__29498\,
            I => \N__29492\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__29495\,
            I => \N__29489\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__29492\,
            I => \N__29486\
        );

    \I__4560\ : Span4Mux_v
    port map (
            O => \N__29489\,
            I => \N__29483\
        );

    \I__4559\ : Span4Mux_h
    port map (
            O => \N__29486\,
            I => \N__29479\
        );

    \I__4558\ : Span4Mux_h
    port map (
            O => \N__29483\,
            I => \N__29476\
        );

    \I__4557\ : InMux
    port map (
            O => \N__29482\,
            I => \N__29473\
        );

    \I__4556\ : Odrv4
    port map (
            O => \N__29479\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__4555\ : Odrv4
    port map (
            O => \N__29476\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__29473\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__4553\ : InMux
    port map (
            O => \N__29466\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__4552\ : InMux
    port map (
            O => \N__29463\,
            I => \N__29460\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__29460\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__4550\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29453\
        );

    \I__4549\ : InMux
    port map (
            O => \N__29456\,
            I => \N__29450\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__29453\,
            I => \N__29447\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__29450\,
            I => \N__29443\
        );

    \I__4546\ : Span4Mux_v
    port map (
            O => \N__29447\,
            I => \N__29440\
        );

    \I__4545\ : InMux
    port map (
            O => \N__29446\,
            I => \N__29437\
        );

    \I__4544\ : Span4Mux_h
    port map (
            O => \N__29443\,
            I => \N__29434\
        );

    \I__4543\ : Span4Mux_v
    port map (
            O => \N__29440\,
            I => \N__29429\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__29437\,
            I => \N__29429\
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__29434\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__4540\ : Odrv4
    port map (
            O => \N__29429\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__4539\ : InMux
    port map (
            O => \N__29424\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__4538\ : InMux
    port map (
            O => \N__29421\,
            I => \N__29418\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__29418\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__4536\ : InMux
    port map (
            O => \N__29415\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__4535\ : InMux
    port map (
            O => \N__29412\,
            I => \N__29409\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__29409\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__4533\ : InMux
    port map (
            O => \N__29406\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__4532\ : InMux
    port map (
            O => \N__29403\,
            I => \N__29400\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__29400\,
            I => \N__29397\
        );

    \I__4530\ : Odrv4
    port map (
            O => \N__29397\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__4529\ : InMux
    port map (
            O => \N__29394\,
            I => \N__29391\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__29391\,
            I => \N__29386\
        );

    \I__4527\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29381\
        );

    \I__4526\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29381\
        );

    \I__4525\ : Odrv4
    port map (
            O => \N__29386\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__29381\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__4523\ : InMux
    port map (
            O => \N__29376\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__4522\ : InMux
    port map (
            O => \N__29373\,
            I => \N__29370\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__29370\,
            I => \N__29367\
        );

    \I__4520\ : Odrv4
    port map (
            O => \N__29367\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__4519\ : InMux
    port map (
            O => \N__29364\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__4518\ : InMux
    port map (
            O => \N__29361\,
            I => \N__29358\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__29358\,
            I => \N__29353\
        );

    \I__4516\ : InMux
    port map (
            O => \N__29357\,
            I => \N__29348\
        );

    \I__4515\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29348\
        );

    \I__4514\ : Span4Mux_v
    port map (
            O => \N__29353\,
            I => \N__29345\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__29348\,
            I => \N__29342\
        );

    \I__4512\ : Odrv4
    port map (
            O => \N__29345\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__4511\ : Odrv12
    port map (
            O => \N__29342\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__4510\ : InMux
    port map (
            O => \N__29337\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__4509\ : CascadeMux
    port map (
            O => \N__29334\,
            I => \N__29331\
        );

    \I__4508\ : InMux
    port map (
            O => \N__29331\,
            I => \N__29326\
        );

    \I__4507\ : InMux
    port map (
            O => \N__29330\,
            I => \N__29323\
        );

    \I__4506\ : InMux
    port map (
            O => \N__29329\,
            I => \N__29320\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__29326\,
            I => \N__29317\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__29323\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__29320\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__4502\ : Odrv4
    port map (
            O => \N__29317\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__4501\ : CascadeMux
    port map (
            O => \N__29310\,
            I => \N__29306\
        );

    \I__4500\ : InMux
    port map (
            O => \N__29309\,
            I => \N__29303\
        );

    \I__4499\ : InMux
    port map (
            O => \N__29306\,
            I => \N__29300\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__29303\,
            I => \N__29296\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__29300\,
            I => \N__29293\
        );

    \I__4496\ : InMux
    port map (
            O => \N__29299\,
            I => \N__29290\
        );

    \I__4495\ : Span4Mux_v
    port map (
            O => \N__29296\,
            I => \N__29283\
        );

    \I__4494\ : Span4Mux_v
    port map (
            O => \N__29293\,
            I => \N__29283\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__29290\,
            I => \N__29283\
        );

    \I__4492\ : Odrv4
    port map (
            O => \N__29283\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__4491\ : InMux
    port map (
            O => \N__29280\,
            I => \N__29277\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__29277\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__4489\ : InMux
    port map (
            O => \N__29274\,
            I => \N__29271\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__29271\,
            I => \N__29267\
        );

    \I__4487\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29264\
        );

    \I__4486\ : Span4Mux_v
    port map (
            O => \N__29267\,
            I => \N__29260\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__29264\,
            I => \N__29257\
        );

    \I__4484\ : InMux
    port map (
            O => \N__29263\,
            I => \N__29254\
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__29260\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__4482\ : Odrv4
    port map (
            O => \N__29257\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__29254\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__4480\ : InMux
    port map (
            O => \N__29247\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__4479\ : InMux
    port map (
            O => \N__29244\,
            I => \N__29241\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__29241\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__4477\ : CascadeMux
    port map (
            O => \N__29238\,
            I => \N__29235\
        );

    \I__4476\ : InMux
    port map (
            O => \N__29235\,
            I => \N__29232\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__29232\,
            I => \N__29228\
        );

    \I__4474\ : InMux
    port map (
            O => \N__29231\,
            I => \N__29225\
        );

    \I__4473\ : Span4Mux_h
    port map (
            O => \N__29228\,
            I => \N__29221\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__29225\,
            I => \N__29218\
        );

    \I__4471\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29215\
        );

    \I__4470\ : Odrv4
    port map (
            O => \N__29221\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__4469\ : Odrv4
    port map (
            O => \N__29218\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__29215\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__4467\ : InMux
    port map (
            O => \N__29208\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__4466\ : InMux
    port map (
            O => \N__29205\,
            I => \N__29202\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__29202\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__29199\,
            I => \N__29196\
        );

    \I__4463\ : InMux
    port map (
            O => \N__29196\,
            I => \N__29193\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__29193\,
            I => \N__29190\
        );

    \I__4461\ : Span4Mux_h
    port map (
            O => \N__29190\,
            I => \N__29186\
        );

    \I__4460\ : InMux
    port map (
            O => \N__29189\,
            I => \N__29182\
        );

    \I__4459\ : Span4Mux_v
    port map (
            O => \N__29186\,
            I => \N__29179\
        );

    \I__4458\ : InMux
    port map (
            O => \N__29185\,
            I => \N__29176\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__29182\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__4456\ : Odrv4
    port map (
            O => \N__29179\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__29176\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__4454\ : InMux
    port map (
            O => \N__29169\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__4453\ : InMux
    port map (
            O => \N__29166\,
            I => \N__29163\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__29163\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__4451\ : CascadeMux
    port map (
            O => \N__29160\,
            I => \N__29156\
        );

    \I__4450\ : InMux
    port map (
            O => \N__29159\,
            I => \N__29153\
        );

    \I__4449\ : InMux
    port map (
            O => \N__29156\,
            I => \N__29150\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__29153\,
            I => \N__29147\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__29150\,
            I => \N__29144\
        );

    \I__4446\ : Span4Mux_v
    port map (
            O => \N__29147\,
            I => \N__29140\
        );

    \I__4445\ : Span4Mux_h
    port map (
            O => \N__29144\,
            I => \N__29137\
        );

    \I__4444\ : InMux
    port map (
            O => \N__29143\,
            I => \N__29134\
        );

    \I__4443\ : Odrv4
    port map (
            O => \N__29140\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__4442\ : Odrv4
    port map (
            O => \N__29137\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__29134\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__4440\ : InMux
    port map (
            O => \N__29127\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__4439\ : InMux
    port map (
            O => \N__29124\,
            I => \N__29121\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__29121\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__4437\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29115\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__29115\,
            I => \N__29110\
        );

    \I__4435\ : InMux
    port map (
            O => \N__29114\,
            I => \N__29105\
        );

    \I__4434\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29105\
        );

    \I__4433\ : Span4Mux_v
    port map (
            O => \N__29110\,
            I => \N__29100\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__29105\,
            I => \N__29100\
        );

    \I__4431\ : Odrv4
    port map (
            O => \N__29100\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__4430\ : InMux
    port map (
            O => \N__29097\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__4429\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29091\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__29091\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__4427\ : InMux
    port map (
            O => \N__29088\,
            I => \N__29084\
        );

    \I__4426\ : CascadeMux
    port map (
            O => \N__29087\,
            I => \N__29080\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__29084\,
            I => \N__29077\
        );

    \I__4424\ : InMux
    port map (
            O => \N__29083\,
            I => \N__29074\
        );

    \I__4423\ : InMux
    port map (
            O => \N__29080\,
            I => \N__29071\
        );

    \I__4422\ : Span4Mux_v
    port map (
            O => \N__29077\,
            I => \N__29066\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__29074\,
            I => \N__29066\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__29071\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__4419\ : Odrv4
    port map (
            O => \N__29066\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__4418\ : InMux
    port map (
            O => \N__29061\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__4417\ : InMux
    port map (
            O => \N__29058\,
            I => \N__29055\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__29055\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__4415\ : InMux
    port map (
            O => \N__29052\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__4414\ : InMux
    port map (
            O => \N__29049\,
            I => \N__29046\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__29046\,
            I => \phase_controller_inst1.stoper_hc.un4_start_0\
        );

    \I__4412\ : InMux
    port map (
            O => \N__29043\,
            I => \N__29034\
        );

    \I__4411\ : InMux
    port map (
            O => \N__29042\,
            I => \N__29034\
        );

    \I__4410\ : InMux
    port map (
            O => \N__29041\,
            I => \N__29034\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__29034\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__4408\ : InMux
    port map (
            O => \N__29031\,
            I => \N__29028\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__29028\,
            I => \N__29025\
        );

    \I__4406\ : Odrv12
    port map (
            O => \N__29025\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__4405\ : CascadeMux
    port map (
            O => \N__29022\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__4404\ : InMux
    port map (
            O => \N__29019\,
            I => \N__29016\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__29016\,
            I => \N__29013\
        );

    \I__4402\ : Span4Mux_v
    port map (
            O => \N__29013\,
            I => \N__29009\
        );

    \I__4401\ : InMux
    port map (
            O => \N__29012\,
            I => \N__29006\
        );

    \I__4400\ : Span4Mux_v
    port map (
            O => \N__29009\,
            I => \N__29001\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__29006\,
            I => \N__29001\
        );

    \I__4398\ : Span4Mux_v
    port map (
            O => \N__29001\,
            I => \N__28998\
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__28998\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__4396\ : InMux
    port map (
            O => \N__28995\,
            I => \N__28992\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__28992\,
            I => \N__28989\
        );

    \I__4394\ : Span4Mux_v
    port map (
            O => \N__28989\,
            I => \N__28985\
        );

    \I__4393\ : InMux
    port map (
            O => \N__28988\,
            I => \N__28982\
        );

    \I__4392\ : Sp12to4
    port map (
            O => \N__28985\,
            I => \N__28978\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__28982\,
            I => \N__28975\
        );

    \I__4390\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28972\
        );

    \I__4389\ : Span12Mux_h
    port map (
            O => \N__28978\,
            I => \N__28967\
        );

    \I__4388\ : Span12Mux_v
    port map (
            O => \N__28975\,
            I => \N__28967\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__28972\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__4386\ : Odrv12
    port map (
            O => \N__28967\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__4385\ : InMux
    port map (
            O => \N__28962\,
            I => \N__28959\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__28959\,
            I => \N__28940\
        );

    \I__4383\ : InMux
    port map (
            O => \N__28958\,
            I => \N__28931\
        );

    \I__4382\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28931\
        );

    \I__4381\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28931\
        );

    \I__4380\ : InMux
    port map (
            O => \N__28955\,
            I => \N__28931\
        );

    \I__4379\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28924\
        );

    \I__4378\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28924\
        );

    \I__4377\ : InMux
    port map (
            O => \N__28952\,
            I => \N__28924\
        );

    \I__4376\ : InMux
    port map (
            O => \N__28951\,
            I => \N__28911\
        );

    \I__4375\ : InMux
    port map (
            O => \N__28950\,
            I => \N__28911\
        );

    \I__4374\ : InMux
    port map (
            O => \N__28949\,
            I => \N__28911\
        );

    \I__4373\ : InMux
    port map (
            O => \N__28948\,
            I => \N__28911\
        );

    \I__4372\ : InMux
    port map (
            O => \N__28947\,
            I => \N__28911\
        );

    \I__4371\ : InMux
    port map (
            O => \N__28946\,
            I => \N__28911\
        );

    \I__4370\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28901\
        );

    \I__4369\ : InMux
    port map (
            O => \N__28944\,
            I => \N__28901\
        );

    \I__4368\ : InMux
    port map (
            O => \N__28943\,
            I => \N__28901\
        );

    \I__4367\ : Span4Mux_h
    port map (
            O => \N__28940\,
            I => \N__28894\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__28931\,
            I => \N__28894\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__28924\,
            I => \N__28894\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__28911\,
            I => \N__28891\
        );

    \I__4363\ : InMux
    port map (
            O => \N__28910\,
            I => \N__28884\
        );

    \I__4362\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28884\
        );

    \I__4361\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28884\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__28901\,
            I => \N__28877\
        );

    \I__4359\ : Span4Mux_v
    port map (
            O => \N__28894\,
            I => \N__28873\
        );

    \I__4358\ : Span4Mux_h
    port map (
            O => \N__28891\,
            I => \N__28868\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__28884\,
            I => \N__28868\
        );

    \I__4356\ : InMux
    port map (
            O => \N__28883\,
            I => \N__28863\
        );

    \I__4355\ : InMux
    port map (
            O => \N__28882\,
            I => \N__28863\
        );

    \I__4354\ : InMux
    port map (
            O => \N__28881\,
            I => \N__28858\
        );

    \I__4353\ : InMux
    port map (
            O => \N__28880\,
            I => \N__28858\
        );

    \I__4352\ : Span4Mux_h
    port map (
            O => \N__28877\,
            I => \N__28855\
        );

    \I__4351\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28852\
        );

    \I__4350\ : Odrv4
    port map (
            O => \N__28873\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__28868\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__28863\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__28858\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__4346\ : Odrv4
    port map (
            O => \N__28855\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__28852\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__4344\ : InMux
    port map (
            O => \N__28839\,
            I => \N__28836\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__28836\,
            I => \N__28833\
        );

    \I__4342\ : Span4Mux_v
    port map (
            O => \N__28833\,
            I => \N__28829\
        );

    \I__4341\ : CascadeMux
    port map (
            O => \N__28832\,
            I => \N__28825\
        );

    \I__4340\ : Span4Mux_v
    port map (
            O => \N__28829\,
            I => \N__28822\
        );

    \I__4339\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28819\
        );

    \I__4338\ : InMux
    port map (
            O => \N__28825\,
            I => \N__28816\
        );

    \I__4337\ : Odrv4
    port map (
            O => \N__28822\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__28819\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__28816\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__4334\ : InMux
    port map (
            O => \N__28809\,
            I => \N__28806\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__28806\,
            I => \N__28803\
        );

    \I__4332\ : Span4Mux_h
    port map (
            O => \N__28803\,
            I => \N__28797\
        );

    \I__4331\ : InMux
    port map (
            O => \N__28802\,
            I => \N__28794\
        );

    \I__4330\ : InMux
    port map (
            O => \N__28801\,
            I => \N__28789\
        );

    \I__4329\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28789\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__28797\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__28794\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__28789\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__28782\,
            I => \N__28779\
        );

    \I__4324\ : InMux
    port map (
            O => \N__28779\,
            I => \N__28773\
        );

    \I__4323\ : InMux
    port map (
            O => \N__28778\,
            I => \N__28770\
        );

    \I__4322\ : InMux
    port map (
            O => \N__28777\,
            I => \N__28767\
        );

    \I__4321\ : InMux
    port map (
            O => \N__28776\,
            I => \N__28762\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__28773\,
            I => \N__28757\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__28770\,
            I => \N__28757\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__28767\,
            I => \N__28754\
        );

    \I__4317\ : InMux
    port map (
            O => \N__28766\,
            I => \N__28751\
        );

    \I__4316\ : InMux
    port map (
            O => \N__28765\,
            I => \N__28748\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__28762\,
            I => \N__28745\
        );

    \I__4314\ : Span4Mux_v
    port map (
            O => \N__28757\,
            I => \N__28740\
        );

    \I__4313\ : Span4Mux_v
    port map (
            O => \N__28754\,
            I => \N__28740\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__28751\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__28748\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__4310\ : Odrv12
    port map (
            O => \N__28745\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__28740\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__4308\ : InMux
    port map (
            O => \N__28731\,
            I => \N__28727\
        );

    \I__4307\ : InMux
    port map (
            O => \N__28730\,
            I => \N__28724\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__28727\,
            I => \N__28721\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__28724\,
            I => \N__28717\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__28721\,
            I => \N__28714\
        );

    \I__4303\ : InMux
    port map (
            O => \N__28720\,
            I => \N__28711\
        );

    \I__4302\ : Odrv12
    port map (
            O => \N__28717\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__28714\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__28711\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__4299\ : InMux
    port map (
            O => \N__28704\,
            I => \N__28700\
        );

    \I__4298\ : CascadeMux
    port map (
            O => \N__28703\,
            I => \N__28697\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__28700\,
            I => \N__28694\
        );

    \I__4296\ : InMux
    port map (
            O => \N__28697\,
            I => \N__28691\
        );

    \I__4295\ : Span4Mux_v
    port map (
            O => \N__28694\,
            I => \N__28688\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__28691\,
            I => \N__28685\
        );

    \I__4293\ : Odrv4
    port map (
            O => \N__28688\,
            I => \phase_controller_inst2.stoper_tr.counter\
        );

    \I__4292\ : Odrv4
    port map (
            O => \N__28685\,
            I => \phase_controller_inst2.stoper_tr.counter\
        );

    \I__4291\ : InMux
    port map (
            O => \N__28680\,
            I => \N__28675\
        );

    \I__4290\ : InMux
    port map (
            O => \N__28679\,
            I => \N__28670\
        );

    \I__4289\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28670\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__28675\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_25\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__28670\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_25\
        );

    \I__4286\ : InMux
    port map (
            O => \N__28665\,
            I => \N__28660\
        );

    \I__4285\ : InMux
    port map (
            O => \N__28664\,
            I => \N__28655\
        );

    \I__4284\ : InMux
    port map (
            O => \N__28663\,
            I => \N__28655\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__28660\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_24\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__28655\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_24\
        );

    \I__4281\ : InMux
    port map (
            O => \N__28650\,
            I => \N__28647\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__28647\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt24\
        );

    \I__4279\ : CascadeMux
    port map (
            O => \N__28644\,
            I => \N__28641\
        );

    \I__4278\ : InMux
    port map (
            O => \N__28641\,
            I => \N__28638\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__28638\,
            I => \N__28635\
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__28635\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt16\
        );

    \I__4275\ : InMux
    port map (
            O => \N__28632\,
            I => \N__28625\
        );

    \I__4274\ : InMux
    port map (
            O => \N__28631\,
            I => \N__28625\
        );

    \I__4273\ : InMux
    port map (
            O => \N__28630\,
            I => \N__28622\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__28625\,
            I => \N__28619\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__28622\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_16\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__28619\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_16\
        );

    \I__4269\ : CascadeMux
    port map (
            O => \N__28614\,
            I => \N__28610\
        );

    \I__4268\ : CascadeMux
    port map (
            O => \N__28613\,
            I => \N__28607\
        );

    \I__4267\ : InMux
    port map (
            O => \N__28610\,
            I => \N__28601\
        );

    \I__4266\ : InMux
    port map (
            O => \N__28607\,
            I => \N__28601\
        );

    \I__4265\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28598\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__28601\,
            I => \N__28595\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__28598\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_17\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__28595\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_17\
        );

    \I__4261\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28587\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__28587\,
            I => \N__28584\
        );

    \I__4259\ : Odrv4
    port map (
            O => \N__28584\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16\
        );

    \I__4258\ : InMux
    port map (
            O => \N__28581\,
            I => \N__28578\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__28578\,
            I => \N__28575\
        );

    \I__4256\ : Span4Mux_h
    port map (
            O => \N__28575\,
            I => \N__28572\
        );

    \I__4255\ : Odrv4
    port map (
            O => \N__28572\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18\
        );

    \I__4254\ : InMux
    port map (
            O => \N__28569\,
            I => \N__28566\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__28566\,
            I => \N__28563\
        );

    \I__4252\ : Odrv12
    port map (
            O => \N__28563\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\
        );

    \I__4251\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28553\
        );

    \I__4250\ : InMux
    port map (
            O => \N__28559\,
            I => \N__28553\
        );

    \I__4249\ : InMux
    port map (
            O => \N__28558\,
            I => \N__28550\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__28553\,
            I => \N__28547\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__28550\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_18\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__28547\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_18\
        );

    \I__4245\ : InMux
    port map (
            O => \N__28542\,
            I => \N__28535\
        );

    \I__4244\ : InMux
    port map (
            O => \N__28541\,
            I => \N__28535\
        );

    \I__4243\ : InMux
    port map (
            O => \N__28540\,
            I => \N__28532\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__28535\,
            I => \N__28529\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__28532\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_19\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__28529\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_19\
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__28524\,
            I => \N__28521\
        );

    \I__4238\ : InMux
    port map (
            O => \N__28521\,
            I => \N__28518\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__28518\,
            I => \N__28515\
        );

    \I__4236\ : Span4Mux_h
    port map (
            O => \N__28515\,
            I => \N__28512\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__28512\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt18\
        );

    \I__4234\ : InMux
    port map (
            O => \N__28509\,
            I => \N__28506\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__28506\,
            I => \N__28503\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__28503\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26\
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__28500\,
            I => \N__28497\
        );

    \I__4230\ : InMux
    port map (
            O => \N__28497\,
            I => \N__28494\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__28494\,
            I => \N__28491\
        );

    \I__4228\ : Span4Mux_h
    port map (
            O => \N__28491\,
            I => \N__28488\
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__28488\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__28485\,
            I => \N__28482\
        );

    \I__4225\ : InMux
    port map (
            O => \N__28482\,
            I => \N__28479\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__28479\,
            I => \N__28476\
        );

    \I__4223\ : Odrv4
    port map (
            O => \N__28476\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30\
        );

    \I__4222\ : InMux
    port map (
            O => \N__28473\,
            I => \bfn_11_10_0_\
        );

    \I__4221\ : InMux
    port map (
            O => \N__28470\,
            I => \N__28465\
        );

    \I__4220\ : InMux
    port map (
            O => \N__28469\,
            I => \N__28462\
        );

    \I__4219\ : InMux
    port map (
            O => \N__28468\,
            I => \N__28459\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__28465\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_31\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__28462\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_31\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__28459\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_31\
        );

    \I__4215\ : InMux
    port map (
            O => \N__28452\,
            I => \N__28447\
        );

    \I__4214\ : InMux
    port map (
            O => \N__28451\,
            I => \N__28444\
        );

    \I__4213\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28441\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__28447\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_30\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__28444\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_30\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__28441\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_30\
        );

    \I__4209\ : InMux
    port map (
            O => \N__28434\,
            I => \N__28431\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__28431\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt30\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__28428\,
            I => \N__28425\
        );

    \I__4206\ : InMux
    port map (
            O => \N__28425\,
            I => \N__28422\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__28422\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24\
        );

    \I__4204\ : InMux
    port map (
            O => \N__28419\,
            I => \N__28413\
        );

    \I__4203\ : InMux
    port map (
            O => \N__28418\,
            I => \N__28408\
        );

    \I__4202\ : InMux
    port map (
            O => \N__28417\,
            I => \N__28408\
        );

    \I__4201\ : InMux
    port map (
            O => \N__28416\,
            I => \N__28405\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__28413\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__28408\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__28405\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28\
        );

    \I__4197\ : InMux
    port map (
            O => \N__28398\,
            I => \N__28393\
        );

    \I__4196\ : InMux
    port map (
            O => \N__28397\,
            I => \N__28390\
        );

    \I__4195\ : InMux
    port map (
            O => \N__28396\,
            I => \N__28387\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__28393\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_29\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__28390\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_29\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__28387\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_29\
        );

    \I__4191\ : InMux
    port map (
            O => \N__28380\,
            I => \N__28375\
        );

    \I__4190\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28372\
        );

    \I__4189\ : InMux
    port map (
            O => \N__28378\,
            I => \N__28369\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__28375\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_28\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__28372\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_28\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__28369\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_28\
        );

    \I__4185\ : InMux
    port map (
            O => \N__28362\,
            I => \N__28359\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__28359\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt28\
        );

    \I__4183\ : InMux
    port map (
            O => \N__28356\,
            I => \N__28352\
        );

    \I__4182\ : InMux
    port map (
            O => \N__28355\,
            I => \N__28349\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__28352\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_11\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__28349\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_11\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__28344\,
            I => \N__28341\
        );

    \I__4178\ : InMux
    port map (
            O => \N__28341\,
            I => \N__28338\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__28338\,
            I => \phase_controller_inst2.stoper_tr.counter_i_11\
        );

    \I__4176\ : InMux
    port map (
            O => \N__28335\,
            I => \N__28331\
        );

    \I__4175\ : InMux
    port map (
            O => \N__28334\,
            I => \N__28328\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__28331\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_12\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__28328\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_12\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__28323\,
            I => \N__28320\
        );

    \I__4171\ : InMux
    port map (
            O => \N__28320\,
            I => \N__28317\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__28317\,
            I => \phase_controller_inst2.stoper_tr.counter_i_12\
        );

    \I__4169\ : InMux
    port map (
            O => \N__28314\,
            I => \N__28310\
        );

    \I__4168\ : InMux
    port map (
            O => \N__28313\,
            I => \N__28307\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__28310\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_13\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__28307\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_13\
        );

    \I__4165\ : CascadeMux
    port map (
            O => \N__28302\,
            I => \N__28299\
        );

    \I__4164\ : InMux
    port map (
            O => \N__28299\,
            I => \N__28296\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__28296\,
            I => \phase_controller_inst2.stoper_tr.counter_i_13\
        );

    \I__4162\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28289\
        );

    \I__4161\ : InMux
    port map (
            O => \N__28292\,
            I => \N__28286\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__28289\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_14\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__28286\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_14\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__28281\,
            I => \N__28278\
        );

    \I__4157\ : InMux
    port map (
            O => \N__28278\,
            I => \N__28275\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__28275\,
            I => \phase_controller_inst2.stoper_tr.counter_i_14\
        );

    \I__4155\ : InMux
    port map (
            O => \N__28272\,
            I => \N__28268\
        );

    \I__4154\ : InMux
    port map (
            O => \N__28271\,
            I => \N__28265\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__28268\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_15\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__28265\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_15\
        );

    \I__4151\ : CascadeMux
    port map (
            O => \N__28260\,
            I => \N__28257\
        );

    \I__4150\ : InMux
    port map (
            O => \N__28257\,
            I => \N__28254\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__28254\,
            I => \phase_controller_inst2.stoper_tr.counter_i_15\
        );

    \I__4148\ : InMux
    port map (
            O => \N__28251\,
            I => \N__28247\
        );

    \I__4147\ : InMux
    port map (
            O => \N__28250\,
            I => \N__28244\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__28247\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_3\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__28244\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_3\
        );

    \I__4144\ : CascadeMux
    port map (
            O => \N__28239\,
            I => \N__28236\
        );

    \I__4143\ : InMux
    port map (
            O => \N__28236\,
            I => \N__28233\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__28233\,
            I => \phase_controller_inst2.stoper_tr.counter_i_3\
        );

    \I__4141\ : InMux
    port map (
            O => \N__28230\,
            I => \N__28226\
        );

    \I__4140\ : InMux
    port map (
            O => \N__28229\,
            I => \N__28223\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__28226\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_4\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__28223\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_4\
        );

    \I__4137\ : CascadeMux
    port map (
            O => \N__28218\,
            I => \N__28215\
        );

    \I__4136\ : InMux
    port map (
            O => \N__28215\,
            I => \N__28212\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__28212\,
            I => \phase_controller_inst2.stoper_tr.counter_i_4\
        );

    \I__4134\ : InMux
    port map (
            O => \N__28209\,
            I => \N__28205\
        );

    \I__4133\ : InMux
    port map (
            O => \N__28208\,
            I => \N__28202\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__28205\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_5\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__28202\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_5\
        );

    \I__4130\ : CascadeMux
    port map (
            O => \N__28197\,
            I => \N__28194\
        );

    \I__4129\ : InMux
    port map (
            O => \N__28194\,
            I => \N__28191\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__28191\,
            I => \phase_controller_inst2.stoper_tr.counter_i_5\
        );

    \I__4127\ : InMux
    port map (
            O => \N__28188\,
            I => \N__28184\
        );

    \I__4126\ : InMux
    port map (
            O => \N__28187\,
            I => \N__28181\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__28184\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_6\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__28181\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_6\
        );

    \I__4123\ : CascadeMux
    port map (
            O => \N__28176\,
            I => \N__28173\
        );

    \I__4122\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28170\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__28170\,
            I => \phase_controller_inst2.stoper_tr.counter_i_6\
        );

    \I__4120\ : InMux
    port map (
            O => \N__28167\,
            I => \N__28163\
        );

    \I__4119\ : InMux
    port map (
            O => \N__28166\,
            I => \N__28160\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__28163\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_7\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__28160\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_7\
        );

    \I__4116\ : CascadeMux
    port map (
            O => \N__28155\,
            I => \N__28152\
        );

    \I__4115\ : InMux
    port map (
            O => \N__28152\,
            I => \N__28149\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__28149\,
            I => \phase_controller_inst2.stoper_tr.counter_i_7\
        );

    \I__4113\ : InMux
    port map (
            O => \N__28146\,
            I => \N__28142\
        );

    \I__4112\ : InMux
    port map (
            O => \N__28145\,
            I => \N__28139\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__28142\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_8\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__28139\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_8\
        );

    \I__4109\ : CascadeMux
    port map (
            O => \N__28134\,
            I => \N__28131\
        );

    \I__4108\ : InMux
    port map (
            O => \N__28131\,
            I => \N__28128\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__28128\,
            I => \phase_controller_inst2.stoper_tr.counter_i_8\
        );

    \I__4106\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28121\
        );

    \I__4105\ : InMux
    port map (
            O => \N__28124\,
            I => \N__28118\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__28121\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_9\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__28118\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_9\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__28113\,
            I => \N__28110\
        );

    \I__4101\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28107\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__28107\,
            I => \phase_controller_inst2.stoper_tr.counter_i_9\
        );

    \I__4099\ : InMux
    port map (
            O => \N__28104\,
            I => \N__28100\
        );

    \I__4098\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28097\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__28100\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_10\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__28097\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_10\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__28092\,
            I => \N__28089\
        );

    \I__4094\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28086\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__28086\,
            I => \phase_controller_inst2.stoper_tr.counter_i_10\
        );

    \I__4092\ : IoInMux
    port map (
            O => \N__28083\,
            I => \N__28080\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__28080\,
            I => \N__28077\
        );

    \I__4090\ : Span4Mux_s1_v
    port map (
            O => \N__28077\,
            I => \N__28074\
        );

    \I__4089\ : Odrv4
    port map (
            O => \N__28074\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__28071\,
            I => \N__28068\
        );

    \I__4087\ : InMux
    port map (
            O => \N__28068\,
            I => \N__28065\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__28065\,
            I => \phase_controller_inst2.stoper_hc.un4_start_0\
        );

    \I__4085\ : InMux
    port map (
            O => \N__28062\,
            I => \N__28056\
        );

    \I__4084\ : InMux
    port map (
            O => \N__28061\,
            I => \N__28056\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__28056\,
            I => \N__28052\
        );

    \I__4082\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28048\
        );

    \I__4081\ : Span4Mux_v
    port map (
            O => \N__28052\,
            I => \N__28045\
        );

    \I__4080\ : InMux
    port map (
            O => \N__28051\,
            I => \N__28042\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__28048\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__28045\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__28042\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__4076\ : InMux
    port map (
            O => \N__28035\,
            I => \N__28030\
        );

    \I__4075\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28024\
        );

    \I__4074\ : InMux
    port map (
            O => \N__28033\,
            I => \N__28021\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__28030\,
            I => \N__28018\
        );

    \I__4072\ : InMux
    port map (
            O => \N__28029\,
            I => \N__28015\
        );

    \I__4071\ : InMux
    port map (
            O => \N__28028\,
            I => \N__28012\
        );

    \I__4070\ : InMux
    port map (
            O => \N__28027\,
            I => \N__28009\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__28024\,
            I => \N__28006\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__28021\,
            I => \N__27999\
        );

    \I__4067\ : Span4Mux_v
    port map (
            O => \N__28018\,
            I => \N__27999\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__28015\,
            I => \N__27999\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__28012\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__28009\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__28006\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__27999\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__4061\ : InMux
    port map (
            O => \N__27990\,
            I => \N__27986\
        );

    \I__4060\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27982\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__27986\,
            I => \N__27979\
        );

    \I__4058\ : InMux
    port map (
            O => \N__27985\,
            I => \N__27976\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__27982\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__27979\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__27976\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__4054\ : InMux
    port map (
            O => \N__27969\,
            I => \N__27965\
        );

    \I__4053\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27962\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__27965\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_0\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__27962\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_0\
        );

    \I__4050\ : CascadeMux
    port map (
            O => \N__27957\,
            I => \N__27954\
        );

    \I__4049\ : InMux
    port map (
            O => \N__27954\,
            I => \N__27951\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__27951\,
            I => \phase_controller_inst2.stoper_tr.counter_i_0\
        );

    \I__4047\ : InMux
    port map (
            O => \N__27948\,
            I => \N__27944\
        );

    \I__4046\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27941\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__27944\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_1\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__27941\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_1\
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__27936\,
            I => \N__27933\
        );

    \I__4042\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27930\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__27930\,
            I => \phase_controller_inst2.stoper_tr.counter_i_1\
        );

    \I__4040\ : InMux
    port map (
            O => \N__27927\,
            I => \N__27923\
        );

    \I__4039\ : InMux
    port map (
            O => \N__27926\,
            I => \N__27920\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__27923\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_2\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__27920\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_2\
        );

    \I__4036\ : CascadeMux
    port map (
            O => \N__27915\,
            I => \N__27912\
        );

    \I__4035\ : InMux
    port map (
            O => \N__27912\,
            I => \N__27909\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__27909\,
            I => \phase_controller_inst2.stoper_tr.counter_i_2\
        );

    \I__4033\ : CascadeMux
    port map (
            O => \N__27906\,
            I => \N__27902\
        );

    \I__4032\ : InMux
    port map (
            O => \N__27905\,
            I => \N__27898\
        );

    \I__4031\ : InMux
    port map (
            O => \N__27902\,
            I => \N__27895\
        );

    \I__4030\ : InMux
    port map (
            O => \N__27901\,
            I => \N__27892\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__27898\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__27895\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__27892\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__4026\ : InMux
    port map (
            O => \N__27885\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__27882\,
            I => \N__27878\
        );

    \I__4024\ : InMux
    port map (
            O => \N__27881\,
            I => \N__27874\
        );

    \I__4023\ : InMux
    port map (
            O => \N__27878\,
            I => \N__27871\
        );

    \I__4022\ : InMux
    port map (
            O => \N__27877\,
            I => \N__27868\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__27874\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__27871\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__27868\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__4018\ : InMux
    port map (
            O => \N__27861\,
            I => \bfn_10_23_0_\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__27858\,
            I => \N__27854\
        );

    \I__4016\ : InMux
    port map (
            O => \N__27857\,
            I => \N__27850\
        );

    \I__4015\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27847\
        );

    \I__4014\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27844\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__27850\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__27847\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__27844\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__4010\ : InMux
    port map (
            O => \N__27837\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__4009\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27830\
        );

    \I__4008\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27827\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__27830\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__27827\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__4005\ : CascadeMux
    port map (
            O => \N__27822\,
            I => \N__27818\
        );

    \I__4004\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27814\
        );

    \I__4003\ : InMux
    port map (
            O => \N__27818\,
            I => \N__27811\
        );

    \I__4002\ : InMux
    port map (
            O => \N__27817\,
            I => \N__27808\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__27814\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__27811\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__27808\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__3998\ : InMux
    port map (
            O => \N__27801\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__3997\ : InMux
    port map (
            O => \N__27798\,
            I => \N__27794\
        );

    \I__3996\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27791\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__27794\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__27791\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__27786\,
            I => \N__27782\
        );

    \I__3992\ : InMux
    port map (
            O => \N__27785\,
            I => \N__27778\
        );

    \I__3991\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27775\
        );

    \I__3990\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27772\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__27778\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__27775\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__27772\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__3986\ : InMux
    port map (
            O => \N__27765\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__3985\ : InMux
    port map (
            O => \N__27762\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__27759\,
            I => \N__27755\
        );

    \I__3983\ : InMux
    port map (
            O => \N__27758\,
            I => \N__27751\
        );

    \I__3982\ : InMux
    port map (
            O => \N__27755\,
            I => \N__27748\
        );

    \I__3981\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27745\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__27751\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__27748\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__27745\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__3977\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27735\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__27735\,
            I => \N__27730\
        );

    \I__3975\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27727\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__27733\,
            I => \N__27724\
        );

    \I__3973\ : Span4Mux_v
    port map (
            O => \N__27730\,
            I => \N__27718\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__27727\,
            I => \N__27718\
        );

    \I__3971\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27713\
        );

    \I__3970\ : InMux
    port map (
            O => \N__27723\,
            I => \N__27713\
        );

    \I__3969\ : Span4Mux_v
    port map (
            O => \N__27718\,
            I => \N__27710\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__27713\,
            I => \N__27707\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__27710\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__3966\ : Odrv12
    port map (
            O => \N__27707\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__3965\ : InMux
    port map (
            O => \N__27702\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__27699\,
            I => \N__27695\
        );

    \I__3963\ : InMux
    port map (
            O => \N__27698\,
            I => \N__27691\
        );

    \I__3962\ : InMux
    port map (
            O => \N__27695\,
            I => \N__27688\
        );

    \I__3961\ : InMux
    port map (
            O => \N__27694\,
            I => \N__27685\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__27691\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__27688\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__27685\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__3957\ : InMux
    port map (
            O => \N__27678\,
            I => \N__27674\
        );

    \I__3956\ : InMux
    port map (
            O => \N__27677\,
            I => \N__27669\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__27674\,
            I => \N__27666\
        );

    \I__3954\ : InMux
    port map (
            O => \N__27673\,
            I => \N__27663\
        );

    \I__3953\ : InMux
    port map (
            O => \N__27672\,
            I => \N__27660\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__27669\,
            I => \N__27657\
        );

    \I__3951\ : Span4Mux_v
    port map (
            O => \N__27666\,
            I => \N__27652\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__27663\,
            I => \N__27652\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__27660\,
            I => \N__27649\
        );

    \I__3948\ : Span4Mux_h
    port map (
            O => \N__27657\,
            I => \N__27646\
        );

    \I__3947\ : Span4Mux_v
    port map (
            O => \N__27652\,
            I => \N__27641\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__27649\,
            I => \N__27641\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__27646\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__27641\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__3943\ : InMux
    port map (
            O => \N__27636\,
            I => \bfn_10_22_0_\
        );

    \I__3942\ : CascadeMux
    port map (
            O => \N__27633\,
            I => \N__27629\
        );

    \I__3941\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27625\
        );

    \I__3940\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27622\
        );

    \I__3939\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27619\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__27625\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__27622\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__27619\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__27612\,
            I => \N__27609\
        );

    \I__3934\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27605\
        );

    \I__3933\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27600\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__27605\,
            I => \N__27597\
        );

    \I__3931\ : InMux
    port map (
            O => \N__27604\,
            I => \N__27594\
        );

    \I__3930\ : InMux
    port map (
            O => \N__27603\,
            I => \N__27591\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__27600\,
            I => \N__27588\
        );

    \I__3928\ : Span4Mux_v
    port map (
            O => \N__27597\,
            I => \N__27581\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__27594\,
            I => \N__27581\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__27591\,
            I => \N__27581\
        );

    \I__3925\ : Span4Mux_v
    port map (
            O => \N__27588\,
            I => \N__27578\
        );

    \I__3924\ : Span4Mux_v
    port map (
            O => \N__27581\,
            I => \N__27575\
        );

    \I__3923\ : Odrv4
    port map (
            O => \N__27578\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__27575\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__3921\ : InMux
    port map (
            O => \N__27570\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__27567\,
            I => \N__27563\
        );

    \I__3919\ : InMux
    port map (
            O => \N__27566\,
            I => \N__27559\
        );

    \I__3918\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27556\
        );

    \I__3917\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27553\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__27559\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__27556\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__27553\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__3913\ : InMux
    port map (
            O => \N__27546\,
            I => \N__27542\
        );

    \I__3912\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27537\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__27542\,
            I => \N__27534\
        );

    \I__3910\ : InMux
    port map (
            O => \N__27541\,
            I => \N__27531\
        );

    \I__3909\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27528\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__27537\,
            I => \N__27523\
        );

    \I__3907\ : Span4Mux_v
    port map (
            O => \N__27534\,
            I => \N__27523\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__27531\,
            I => \N__27518\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__27528\,
            I => \N__27518\
        );

    \I__3904\ : Odrv4
    port map (
            O => \N__27523\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__3903\ : Odrv12
    port map (
            O => \N__27518\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__3902\ : InMux
    port map (
            O => \N__27513\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__27510\,
            I => \N__27506\
        );

    \I__3900\ : InMux
    port map (
            O => \N__27509\,
            I => \N__27502\
        );

    \I__3899\ : InMux
    port map (
            O => \N__27506\,
            I => \N__27499\
        );

    \I__3898\ : InMux
    port map (
            O => \N__27505\,
            I => \N__27496\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__27502\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__27499\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__27496\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__27489\,
            I => \N__27486\
        );

    \I__3893\ : InMux
    port map (
            O => \N__27486\,
            I => \N__27483\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__27483\,
            I => \N__27478\
        );

    \I__3891\ : InMux
    port map (
            O => \N__27482\,
            I => \N__27475\
        );

    \I__3890\ : InMux
    port map (
            O => \N__27481\,
            I => \N__27471\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__27478\,
            I => \N__27466\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__27475\,
            I => \N__27466\
        );

    \I__3887\ : InMux
    port map (
            O => \N__27474\,
            I => \N__27463\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__27471\,
            I => \N__27460\
        );

    \I__3885\ : Sp12to4
    port map (
            O => \N__27466\,
            I => \N__27455\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__27463\,
            I => \N__27455\
        );

    \I__3883\ : Odrv4
    port map (
            O => \N__27460\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__3882\ : Odrv12
    port map (
            O => \N__27455\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__3881\ : InMux
    port map (
            O => \N__27450\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__27447\,
            I => \N__27443\
        );

    \I__3879\ : InMux
    port map (
            O => \N__27446\,
            I => \N__27439\
        );

    \I__3878\ : InMux
    port map (
            O => \N__27443\,
            I => \N__27436\
        );

    \I__3877\ : InMux
    port map (
            O => \N__27442\,
            I => \N__27433\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__27439\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__27436\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__27433\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__3873\ : InMux
    port map (
            O => \N__27426\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__3872\ : CascadeMux
    port map (
            O => \N__27423\,
            I => \N__27419\
        );

    \I__3871\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27415\
        );

    \I__3870\ : InMux
    port map (
            O => \N__27419\,
            I => \N__27412\
        );

    \I__3869\ : InMux
    port map (
            O => \N__27418\,
            I => \N__27409\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__27415\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__27412\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__27409\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__3865\ : InMux
    port map (
            O => \N__27402\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__27399\,
            I => \N__27395\
        );

    \I__3863\ : InMux
    port map (
            O => \N__27398\,
            I => \N__27391\
        );

    \I__3862\ : InMux
    port map (
            O => \N__27395\,
            I => \N__27388\
        );

    \I__3861\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27385\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__27391\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__27388\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__27385\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__3857\ : InMux
    port map (
            O => \N__27378\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__3856\ : CascadeMux
    port map (
            O => \N__27375\,
            I => \N__27371\
        );

    \I__3855\ : InMux
    port map (
            O => \N__27374\,
            I => \N__27367\
        );

    \I__3854\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27364\
        );

    \I__3853\ : InMux
    port map (
            O => \N__27370\,
            I => \N__27361\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__27367\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__27364\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__27361\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__3849\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27350\
        );

    \I__3848\ : CascadeMux
    port map (
            O => \N__27353\,
            I => \N__27347\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__27350\,
            I => \N__27343\
        );

    \I__3846\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27340\
        );

    \I__3845\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27337\
        );

    \I__3844\ : Span4Mux_v
    port map (
            O => \N__27343\,
            I => \N__27330\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__27340\,
            I => \N__27330\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__27337\,
            I => \N__27330\
        );

    \I__3841\ : Span4Mux_v
    port map (
            O => \N__27330\,
            I => \N__27326\
        );

    \I__3840\ : InMux
    port map (
            O => \N__27329\,
            I => \N__27323\
        );

    \I__3839\ : Odrv4
    port map (
            O => \N__27326\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__27323\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__3837\ : InMux
    port map (
            O => \N__27318\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__27315\,
            I => \N__27311\
        );

    \I__3835\ : InMux
    port map (
            O => \N__27314\,
            I => \N__27307\
        );

    \I__3834\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27304\
        );

    \I__3833\ : InMux
    port map (
            O => \N__27310\,
            I => \N__27301\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__27307\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__27304\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__27301\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__27294\,
            I => \N__27290\
        );

    \I__3828\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27286\
        );

    \I__3827\ : InMux
    port map (
            O => \N__27290\,
            I => \N__27283\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__27289\,
            I => \N__27280\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__27286\,
            I => \N__27276\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__27283\,
            I => \N__27273\
        );

    \I__3823\ : InMux
    port map (
            O => \N__27280\,
            I => \N__27270\
        );

    \I__3822\ : InMux
    port map (
            O => \N__27279\,
            I => \N__27267\
        );

    \I__3821\ : Span4Mux_v
    port map (
            O => \N__27276\,
            I => \N__27264\
        );

    \I__3820\ : Sp12to4
    port map (
            O => \N__27273\,
            I => \N__27257\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__27270\,
            I => \N__27257\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__27267\,
            I => \N__27257\
        );

    \I__3817\ : Odrv4
    port map (
            O => \N__27264\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__3816\ : Odrv12
    port map (
            O => \N__27257\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__3815\ : InMux
    port map (
            O => \N__27252\,
            I => \bfn_10_21_0_\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__27249\,
            I => \N__27245\
        );

    \I__3813\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27241\
        );

    \I__3812\ : InMux
    port map (
            O => \N__27245\,
            I => \N__27238\
        );

    \I__3811\ : InMux
    port map (
            O => \N__27244\,
            I => \N__27235\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__27241\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__27238\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__27235\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__27228\,
            I => \N__27223\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__27227\,
            I => \N__27220\
        );

    \I__3805\ : InMux
    port map (
            O => \N__27226\,
            I => \N__27217\
        );

    \I__3804\ : InMux
    port map (
            O => \N__27223\,
            I => \N__27214\
        );

    \I__3803\ : InMux
    port map (
            O => \N__27220\,
            I => \N__27210\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__27217\,
            I => \N__27207\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__27214\,
            I => \N__27204\
        );

    \I__3800\ : InMux
    port map (
            O => \N__27213\,
            I => \N__27201\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__27210\,
            I => \N__27198\
        );

    \I__3798\ : Span4Mux_v
    port map (
            O => \N__27207\,
            I => \N__27195\
        );

    \I__3797\ : Sp12to4
    port map (
            O => \N__27204\,
            I => \N__27190\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__27201\,
            I => \N__27190\
        );

    \I__3795\ : Odrv12
    port map (
            O => \N__27198\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__3794\ : Odrv4
    port map (
            O => \N__27195\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__3793\ : Odrv12
    port map (
            O => \N__27190\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__3792\ : InMux
    port map (
            O => \N__27183\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__3791\ : CascadeMux
    port map (
            O => \N__27180\,
            I => \N__27176\
        );

    \I__3790\ : InMux
    port map (
            O => \N__27179\,
            I => \N__27172\
        );

    \I__3789\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27169\
        );

    \I__3788\ : InMux
    port map (
            O => \N__27175\,
            I => \N__27166\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__27172\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__27169\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__27166\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__3784\ : InMux
    port map (
            O => \N__27159\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__27156\,
            I => \N__27152\
        );

    \I__3782\ : InMux
    port map (
            O => \N__27155\,
            I => \N__27148\
        );

    \I__3781\ : InMux
    port map (
            O => \N__27152\,
            I => \N__27145\
        );

    \I__3780\ : InMux
    port map (
            O => \N__27151\,
            I => \N__27142\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__27148\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__27145\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__27142\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__3776\ : InMux
    port map (
            O => \N__27135\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__3775\ : CascadeMux
    port map (
            O => \N__27132\,
            I => \N__27128\
        );

    \I__3774\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27124\
        );

    \I__3773\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27121\
        );

    \I__3772\ : InMux
    port map (
            O => \N__27127\,
            I => \N__27118\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__27124\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__27121\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__27118\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__27111\,
            I => \N__27107\
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__27110\,
            I => \N__27104\
        );

    \I__3766\ : InMux
    port map (
            O => \N__27107\,
            I => \N__27100\
        );

    \I__3765\ : InMux
    port map (
            O => \N__27104\,
            I => \N__27095\
        );

    \I__3764\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27095\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__27100\,
            I => \N__27089\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__27095\,
            I => \N__27089\
        );

    \I__3761\ : InMux
    port map (
            O => \N__27094\,
            I => \N__27086\
        );

    \I__3760\ : Span4Mux_v
    port map (
            O => \N__27089\,
            I => \N__27081\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__27086\,
            I => \N__27081\
        );

    \I__3758\ : Odrv4
    port map (
            O => \N__27081\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__3757\ : InMux
    port map (
            O => \N__27078\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__27075\,
            I => \N__27071\
        );

    \I__3755\ : InMux
    port map (
            O => \N__27074\,
            I => \N__27067\
        );

    \I__3754\ : InMux
    port map (
            O => \N__27071\,
            I => \N__27064\
        );

    \I__3753\ : InMux
    port map (
            O => \N__27070\,
            I => \N__27061\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__27067\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__27064\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__27061\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__3749\ : InMux
    port map (
            O => \N__27054\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__27051\,
            I => \N__27047\
        );

    \I__3747\ : InMux
    port map (
            O => \N__27050\,
            I => \N__27043\
        );

    \I__3746\ : InMux
    port map (
            O => \N__27047\,
            I => \N__27040\
        );

    \I__3745\ : InMux
    port map (
            O => \N__27046\,
            I => \N__27037\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__27043\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__27040\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__27037\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__3741\ : InMux
    port map (
            O => \N__27030\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__3740\ : InMux
    port map (
            O => \N__27027\,
            I => \N__27024\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__27024\,
            I => \N__27021\
        );

    \I__3738\ : Span4Mux_h
    port map (
            O => \N__27021\,
            I => \N__27018\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__27018\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__3736\ : CascadeMux
    port map (
            O => \N__27015\,
            I => \N__27011\
        );

    \I__3735\ : InMux
    port map (
            O => \N__27014\,
            I => \N__27008\
        );

    \I__3734\ : InMux
    port map (
            O => \N__27011\,
            I => \N__27003\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__27008\,
            I => \N__27000\
        );

    \I__3732\ : InMux
    port map (
            O => \N__27007\,
            I => \N__26997\
        );

    \I__3731\ : InMux
    port map (
            O => \N__27006\,
            I => \N__26994\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__27003\,
            I => \N__26991\
        );

    \I__3729\ : Span4Mux_v
    port map (
            O => \N__27000\,
            I => \N__26988\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__26997\,
            I => \N__26983\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__26994\,
            I => \N__26983\
        );

    \I__3726\ : Odrv4
    port map (
            O => \N__26991\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__3725\ : Odrv4
    port map (
            O => \N__26988\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__3724\ : Odrv12
    port map (
            O => \N__26983\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__3723\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26973\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__26973\,
            I => \N__26969\
        );

    \I__3721\ : InMux
    port map (
            O => \N__26972\,
            I => \N__26966\
        );

    \I__3720\ : Span4Mux_v
    port map (
            O => \N__26969\,
            I => \N__26959\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__26966\,
            I => \N__26959\
        );

    \I__3718\ : InMux
    port map (
            O => \N__26965\,
            I => \N__26954\
        );

    \I__3717\ : InMux
    port map (
            O => \N__26964\,
            I => \N__26954\
        );

    \I__3716\ : Span4Mux_v
    port map (
            O => \N__26959\,
            I => \N__26951\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__26954\,
            I => \N__26948\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__26951\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__3713\ : Odrv12
    port map (
            O => \N__26948\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__3712\ : InMux
    port map (
            O => \N__26943\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__26940\,
            I => \N__26936\
        );

    \I__3710\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26932\
        );

    \I__3709\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26929\
        );

    \I__3708\ : InMux
    port map (
            O => \N__26935\,
            I => \N__26926\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__26932\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__26929\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__26926\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__3704\ : InMux
    port map (
            O => \N__26919\,
            I => \N__26913\
        );

    \I__3703\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26910\
        );

    \I__3702\ : InMux
    port map (
            O => \N__26917\,
            I => \N__26907\
        );

    \I__3701\ : InMux
    port map (
            O => \N__26916\,
            I => \N__26904\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__26913\,
            I => \N__26901\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__26910\,
            I => \N__26894\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__26907\,
            I => \N__26894\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__26904\,
            I => \N__26894\
        );

    \I__3696\ : Odrv4
    port map (
            O => \N__26901\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__3695\ : Odrv12
    port map (
            O => \N__26894\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__3694\ : InMux
    port map (
            O => \N__26889\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__3693\ : CascadeMux
    port map (
            O => \N__26886\,
            I => \N__26882\
        );

    \I__3692\ : InMux
    port map (
            O => \N__26885\,
            I => \N__26878\
        );

    \I__3691\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26875\
        );

    \I__3690\ : InMux
    port map (
            O => \N__26881\,
            I => \N__26872\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__26878\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__26875\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__26872\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__3686\ : CascadeMux
    port map (
            O => \N__26865\,
            I => \N__26862\
        );

    \I__3685\ : InMux
    port map (
            O => \N__26862\,
            I => \N__26858\
        );

    \I__3684\ : InMux
    port map (
            O => \N__26861\,
            I => \N__26853\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__26858\,
            I => \N__26850\
        );

    \I__3682\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26847\
        );

    \I__3681\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26844\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__26853\,
            I => \N__26841\
        );

    \I__3679\ : Sp12to4
    port map (
            O => \N__26850\,
            I => \N__26834\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__26847\,
            I => \N__26834\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__26844\,
            I => \N__26834\
        );

    \I__3676\ : Odrv4
    port map (
            O => \N__26841\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__3675\ : Odrv12
    port map (
            O => \N__26834\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__3674\ : InMux
    port map (
            O => \N__26829\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__26826\,
            I => \N__26822\
        );

    \I__3672\ : InMux
    port map (
            O => \N__26825\,
            I => \N__26818\
        );

    \I__3671\ : InMux
    port map (
            O => \N__26822\,
            I => \N__26815\
        );

    \I__3670\ : InMux
    port map (
            O => \N__26821\,
            I => \N__26812\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__26818\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__26815\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__26812\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__3666\ : CascadeMux
    port map (
            O => \N__26805\,
            I => \N__26800\
        );

    \I__3665\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26796\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__26803\,
            I => \N__26793\
        );

    \I__3663\ : InMux
    port map (
            O => \N__26800\,
            I => \N__26788\
        );

    \I__3662\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26788\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__26796\,
            I => \N__26785\
        );

    \I__3660\ : InMux
    port map (
            O => \N__26793\,
            I => \N__26782\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__26788\,
            I => \N__26779\
        );

    \I__3658\ : Span4Mux_v
    port map (
            O => \N__26785\,
            I => \N__26776\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__26782\,
            I => \N__26771\
        );

    \I__3656\ : Span4Mux_v
    port map (
            O => \N__26779\,
            I => \N__26771\
        );

    \I__3655\ : Span4Mux_v
    port map (
            O => \N__26776\,
            I => \N__26768\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__26771\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__26768\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__3652\ : InMux
    port map (
            O => \N__26763\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__3651\ : CascadeMux
    port map (
            O => \N__26760\,
            I => \N__26756\
        );

    \I__3650\ : InMux
    port map (
            O => \N__26759\,
            I => \N__26752\
        );

    \I__3649\ : InMux
    port map (
            O => \N__26756\,
            I => \N__26749\
        );

    \I__3648\ : InMux
    port map (
            O => \N__26755\,
            I => \N__26746\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__26752\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__26749\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__26746\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__3644\ : CascadeMux
    port map (
            O => \N__26739\,
            I => \N__26736\
        );

    \I__3643\ : InMux
    port map (
            O => \N__26736\,
            I => \N__26731\
        );

    \I__3642\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26727\
        );

    \I__3641\ : InMux
    port map (
            O => \N__26734\,
            I => \N__26724\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__26731\,
            I => \N__26721\
        );

    \I__3639\ : InMux
    port map (
            O => \N__26730\,
            I => \N__26718\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__26727\,
            I => \N__26713\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__26724\,
            I => \N__26713\
        );

    \I__3636\ : Span4Mux_v
    port map (
            O => \N__26721\,
            I => \N__26706\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__26718\,
            I => \N__26706\
        );

    \I__3634\ : Span4Mux_h
    port map (
            O => \N__26713\,
            I => \N__26706\
        );

    \I__3633\ : Span4Mux_v
    port map (
            O => \N__26706\,
            I => \N__26703\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__26703\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__3631\ : InMux
    port map (
            O => \N__26700\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__3630\ : CascadeMux
    port map (
            O => \N__26697\,
            I => \N__26693\
        );

    \I__3629\ : InMux
    port map (
            O => \N__26696\,
            I => \N__26689\
        );

    \I__3628\ : InMux
    port map (
            O => \N__26693\,
            I => \N__26686\
        );

    \I__3627\ : InMux
    port map (
            O => \N__26692\,
            I => \N__26683\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__26689\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__26686\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__26683\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__3623\ : InMux
    port map (
            O => \N__26676\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__26673\,
            I => \N__26670\
        );

    \I__3621\ : InMux
    port map (
            O => \N__26670\,
            I => \N__26667\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__26667\,
            I => \N__26664\
        );

    \I__3619\ : Odrv12
    port map (
            O => \N__26664\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__3618\ : InMux
    port map (
            O => \N__26661\,
            I => \N__26658\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__26658\,
            I => \N__26655\
        );

    \I__3616\ : Odrv4
    port map (
            O => \N__26655\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__3615\ : InMux
    port map (
            O => \N__26652\,
            I => \N__26649\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__26649\,
            I => \N__26646\
        );

    \I__3613\ : Span4Mux_v
    port map (
            O => \N__26646\,
            I => \N__26643\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__26643\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__26640\,
            I => \N__26637\
        );

    \I__3610\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26634\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__26634\,
            I => \N__26631\
        );

    \I__3608\ : Span4Mux_h
    port map (
            O => \N__26631\,
            I => \N__26628\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__26628\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__26625\,
            I => \N__26622\
        );

    \I__3605\ : InMux
    port map (
            O => \N__26622\,
            I => \N__26619\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__26619\,
            I => \N__26616\
        );

    \I__3603\ : Span4Mux_v
    port map (
            O => \N__26616\,
            I => \N__26613\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__26613\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__3601\ : CascadeMux
    port map (
            O => \N__26610\,
            I => \N__26607\
        );

    \I__3600\ : InMux
    port map (
            O => \N__26607\,
            I => \N__26604\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__26604\,
            I => \N__26601\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__26601\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\
        );

    \I__3597\ : CascadeMux
    port map (
            O => \N__26598\,
            I => \N__26595\
        );

    \I__3596\ : InMux
    port map (
            O => \N__26595\,
            I => \N__26592\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__26592\,
            I => \N__26589\
        );

    \I__3594\ : Span4Mux_h
    port map (
            O => \N__26589\,
            I => \N__26586\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__26586\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__26583\,
            I => \N__26580\
        );

    \I__3591\ : InMux
    port map (
            O => \N__26580\,
            I => \N__26577\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__26577\,
            I => \N__26574\
        );

    \I__3589\ : Span4Mux_h
    port map (
            O => \N__26574\,
            I => \N__26571\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__26571\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__26568\,
            I => \N__26565\
        );

    \I__3586\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26562\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__26562\,
            I => \N__26559\
        );

    \I__3584\ : Odrv4
    port map (
            O => \N__26559\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__3583\ : InMux
    port map (
            O => \N__26556\,
            I => \N__26553\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__26553\,
            I => \N__26550\
        );

    \I__3581\ : Span4Mux_h
    port map (
            O => \N__26550\,
            I => \N__26547\
        );

    \I__3580\ : Odrv4
    port map (
            O => \N__26547\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\
        );

    \I__3579\ : InMux
    port map (
            O => \N__26544\,
            I => \N__26541\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__26541\,
            I => \N__26538\
        );

    \I__3577\ : Span4Mux_v
    port map (
            O => \N__26538\,
            I => \N__26535\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__26535\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__26532\,
            I => \N__26529\
        );

    \I__3574\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26526\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__26526\,
            I => \N__26523\
        );

    \I__3572\ : Odrv12
    port map (
            O => \N__26523\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__26520\,
            I => \N__26517\
        );

    \I__3570\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26514\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__26514\,
            I => \N__26511\
        );

    \I__3568\ : Span4Mux_h
    port map (
            O => \N__26511\,
            I => \N__26508\
        );

    \I__3567\ : Span4Mux_h
    port map (
            O => \N__26508\,
            I => \N__26505\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__26505\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__3565\ : CascadeMux
    port map (
            O => \N__26502\,
            I => \N__26499\
        );

    \I__3564\ : InMux
    port map (
            O => \N__26499\,
            I => \N__26496\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__26496\,
            I => \N__26493\
        );

    \I__3562\ : Odrv4
    port map (
            O => \N__26493\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__26490\,
            I => \N__26487\
        );

    \I__3560\ : InMux
    port map (
            O => \N__26487\,
            I => \N__26484\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__26484\,
            I => \N__26481\
        );

    \I__3558\ : Odrv4
    port map (
            O => \N__26481\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__3557\ : CascadeMux
    port map (
            O => \N__26478\,
            I => \N__26475\
        );

    \I__3556\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26472\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__26472\,
            I => \N__26469\
        );

    \I__3554\ : Span4Mux_h
    port map (
            O => \N__26469\,
            I => \N__26466\
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__26466\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__26463\,
            I => \N__26460\
        );

    \I__3551\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26457\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__26457\,
            I => \N__26454\
        );

    \I__3549\ : Span4Mux_h
    port map (
            O => \N__26454\,
            I => \N__26451\
        );

    \I__3548\ : Odrv4
    port map (
            O => \N__26451\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__26448\,
            I => \N__26445\
        );

    \I__3546\ : InMux
    port map (
            O => \N__26445\,
            I => \N__26442\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__26442\,
            I => \N__26439\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__26439\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__26436\,
            I => \N__26433\
        );

    \I__3542\ : InMux
    port map (
            O => \N__26433\,
            I => \N__26430\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__26430\,
            I => \N__26427\
        );

    \I__3540\ : Odrv4
    port map (
            O => \N__26427\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__3539\ : CascadeMux
    port map (
            O => \N__26424\,
            I => \N__26421\
        );

    \I__3538\ : InMux
    port map (
            O => \N__26421\,
            I => \N__26418\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__26418\,
            I => \N__26415\
        );

    \I__3536\ : Span4Mux_v
    port map (
            O => \N__26415\,
            I => \N__26412\
        );

    \I__3535\ : Odrv4
    port map (
            O => \N__26412\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__3534\ : InMux
    port map (
            O => \N__26409\,
            I => \N__26406\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__26406\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__3532\ : CascadeMux
    port map (
            O => \N__26403\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__3531\ : InMux
    port map (
            O => \N__26400\,
            I => \N__26396\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__26399\,
            I => \N__26393\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__26396\,
            I => \N__26390\
        );

    \I__3528\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26387\
        );

    \I__3527\ : Span4Mux_v
    port map (
            O => \N__26390\,
            I => \N__26382\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__26387\,
            I => \N__26382\
        );

    \I__3525\ : Span4Mux_v
    port map (
            O => \N__26382\,
            I => \N__26379\
        );

    \I__3524\ : Span4Mux_v
    port map (
            O => \N__26379\,
            I => \N__26376\
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__26376\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__3522\ : InMux
    port map (
            O => \N__26373\,
            I => \N__26370\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__26370\,
            I => \N__26367\
        );

    \I__3520\ : Span4Mux_h
    port map (
            O => \N__26367\,
            I => \N__26364\
        );

    \I__3519\ : Span4Mux_v
    port map (
            O => \N__26364\,
            I => \N__26361\
        );

    \I__3518\ : Odrv4
    port map (
            O => \N__26361\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__26358\,
            I => \N__26355\
        );

    \I__3516\ : InMux
    port map (
            O => \N__26355\,
            I => \N__26352\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__26352\,
            I => \N__26349\
        );

    \I__3514\ : Span4Mux_h
    port map (
            O => \N__26349\,
            I => \N__26346\
        );

    \I__3513\ : Span4Mux_h
    port map (
            O => \N__26346\,
            I => \N__26343\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__26343\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__26340\,
            I => \N__26337\
        );

    \I__3510\ : InMux
    port map (
            O => \N__26337\,
            I => \N__26334\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__26334\,
            I => \N__26331\
        );

    \I__3508\ : Span4Mux_v
    port map (
            O => \N__26331\,
            I => \N__26328\
        );

    \I__3507\ : Odrv4
    port map (
            O => \N__26328\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\
        );

    \I__3506\ : InMux
    port map (
            O => \N__26325\,
            I => \N__26322\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__26322\,
            I => \N__26319\
        );

    \I__3504\ : Odrv4
    port map (
            O => \N__26319\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__26316\,
            I => \N__26313\
        );

    \I__3502\ : InMux
    port map (
            O => \N__26313\,
            I => \N__26310\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__26310\,
            I => \N__26307\
        );

    \I__3500\ : Span4Mux_h
    port map (
            O => \N__26307\,
            I => \N__26304\
        );

    \I__3499\ : Odrv4
    port map (
            O => \N__26304\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\
        );

    \I__3498\ : InMux
    port map (
            O => \N__26301\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_28\
        );

    \I__3497\ : InMux
    port map (
            O => \N__26298\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_29\
        );

    \I__3496\ : InMux
    port map (
            O => \N__26295\,
            I => \N__26255\
        );

    \I__3495\ : InMux
    port map (
            O => \N__26294\,
            I => \N__26255\
        );

    \I__3494\ : InMux
    port map (
            O => \N__26293\,
            I => \N__26255\
        );

    \I__3493\ : InMux
    port map (
            O => \N__26292\,
            I => \N__26255\
        );

    \I__3492\ : InMux
    port map (
            O => \N__26291\,
            I => \N__26246\
        );

    \I__3491\ : InMux
    port map (
            O => \N__26290\,
            I => \N__26246\
        );

    \I__3490\ : InMux
    port map (
            O => \N__26289\,
            I => \N__26246\
        );

    \I__3489\ : InMux
    port map (
            O => \N__26288\,
            I => \N__26246\
        );

    \I__3488\ : InMux
    port map (
            O => \N__26287\,
            I => \N__26237\
        );

    \I__3487\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26237\
        );

    \I__3486\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26237\
        );

    \I__3485\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26237\
        );

    \I__3484\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26228\
        );

    \I__3483\ : InMux
    port map (
            O => \N__26282\,
            I => \N__26228\
        );

    \I__3482\ : InMux
    port map (
            O => \N__26281\,
            I => \N__26228\
        );

    \I__3481\ : InMux
    port map (
            O => \N__26280\,
            I => \N__26228\
        );

    \I__3480\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26219\
        );

    \I__3479\ : InMux
    port map (
            O => \N__26278\,
            I => \N__26219\
        );

    \I__3478\ : InMux
    port map (
            O => \N__26277\,
            I => \N__26219\
        );

    \I__3477\ : InMux
    port map (
            O => \N__26276\,
            I => \N__26219\
        );

    \I__3476\ : InMux
    port map (
            O => \N__26275\,
            I => \N__26210\
        );

    \I__3475\ : InMux
    port map (
            O => \N__26274\,
            I => \N__26210\
        );

    \I__3474\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26210\
        );

    \I__3473\ : InMux
    port map (
            O => \N__26272\,
            I => \N__26210\
        );

    \I__3472\ : InMux
    port map (
            O => \N__26271\,
            I => \N__26201\
        );

    \I__3471\ : InMux
    port map (
            O => \N__26270\,
            I => \N__26201\
        );

    \I__3470\ : InMux
    port map (
            O => \N__26269\,
            I => \N__26201\
        );

    \I__3469\ : InMux
    port map (
            O => \N__26268\,
            I => \N__26201\
        );

    \I__3468\ : InMux
    port map (
            O => \N__26267\,
            I => \N__26192\
        );

    \I__3467\ : InMux
    port map (
            O => \N__26266\,
            I => \N__26192\
        );

    \I__3466\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26192\
        );

    \I__3465\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26192\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__26255\,
            I => \N__26183\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__26246\,
            I => \N__26183\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__26237\,
            I => \N__26183\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__26228\,
            I => \N__26183\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__26219\,
            I => \phase_controller_inst2.stoper_tr.start_latched_i_0\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__26210\,
            I => \phase_controller_inst2.stoper_tr.start_latched_i_0\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__26201\,
            I => \phase_controller_inst2.stoper_tr.start_latched_i_0\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__26192\,
            I => \phase_controller_inst2.stoper_tr.start_latched_i_0\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__26183\,
            I => \phase_controller_inst2.stoper_tr.start_latched_i_0\
        );

    \I__3455\ : InMux
    port map (
            O => \N__26172\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_30\
        );

    \I__3454\ : CEMux
    port map (
            O => \N__26169\,
            I => \N__26157\
        );

    \I__3453\ : CEMux
    port map (
            O => \N__26168\,
            I => \N__26157\
        );

    \I__3452\ : CEMux
    port map (
            O => \N__26167\,
            I => \N__26157\
        );

    \I__3451\ : CEMux
    port map (
            O => \N__26166\,
            I => \N__26157\
        );

    \I__3450\ : GlobalMux
    port map (
            O => \N__26157\,
            I => \N__26154\
        );

    \I__3449\ : gio2CtrlBuf
    port map (
            O => \N__26154\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0_g\
        );

    \I__3448\ : InMux
    port map (
            O => \N__26151\,
            I => \N__26147\
        );

    \I__3447\ : InMux
    port map (
            O => \N__26150\,
            I => \N__26144\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__26147\,
            I => \N__26141\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__26144\,
            I => \N__26138\
        );

    \I__3444\ : Span4Mux_v
    port map (
            O => \N__26141\,
            I => \N__26135\
        );

    \I__3443\ : Span4Mux_v
    port map (
            O => \N__26138\,
            I => \N__26132\
        );

    \I__3442\ : Span4Mux_h
    port map (
            O => \N__26135\,
            I => \N__26129\
        );

    \I__3441\ : Span4Mux_h
    port map (
            O => \N__26132\,
            I => \N__26126\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__26129\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__3439\ : Odrv4
    port map (
            O => \N__26126\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__3438\ : InMux
    port map (
            O => \N__26121\,
            I => \N__26118\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__26118\,
            I => \N__26114\
        );

    \I__3436\ : InMux
    port map (
            O => \N__26117\,
            I => \N__26111\
        );

    \I__3435\ : Sp12to4
    port map (
            O => \N__26114\,
            I => \N__26106\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__26111\,
            I => \N__26106\
        );

    \I__3433\ : Odrv12
    port map (
            O => \N__26106\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__3432\ : InMux
    port map (
            O => \N__26103\,
            I => \N__26099\
        );

    \I__3431\ : InMux
    port map (
            O => \N__26102\,
            I => \N__26096\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__26099\,
            I => \N__26093\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__26096\,
            I => \N__26090\
        );

    \I__3428\ : Span12Mux_s5_h
    port map (
            O => \N__26093\,
            I => \N__26087\
        );

    \I__3427\ : Odrv12
    port map (
            O => \N__26090\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__3426\ : Odrv12
    port map (
            O => \N__26087\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__3425\ : InMux
    port map (
            O => \N__26082\,
            I => \N__26078\
        );

    \I__3424\ : InMux
    port map (
            O => \N__26081\,
            I => \N__26075\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__26078\,
            I => \N__26072\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__26075\,
            I => \N__26069\
        );

    \I__3421\ : Span4Mux_s3_h
    port map (
            O => \N__26072\,
            I => \N__26066\
        );

    \I__3420\ : Odrv12
    port map (
            O => \N__26069\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__3419\ : Odrv4
    port map (
            O => \N__26066\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__3418\ : InMux
    port map (
            O => \N__26061\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_19\
        );

    \I__3417\ : InMux
    port map (
            O => \N__26058\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_20\
        );

    \I__3416\ : InMux
    port map (
            O => \N__26055\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_21\
        );

    \I__3415\ : InMux
    port map (
            O => \N__26052\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_22\
        );

    \I__3414\ : InMux
    port map (
            O => \N__26049\,
            I => \bfn_10_10_0_\
        );

    \I__3413\ : InMux
    port map (
            O => \N__26046\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_24\
        );

    \I__3412\ : InMux
    port map (
            O => \N__26043\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_25\
        );

    \I__3411\ : InMux
    port map (
            O => \N__26040\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_26\
        );

    \I__3410\ : InMux
    port map (
            O => \N__26037\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_27\
        );

    \I__3409\ : InMux
    port map (
            O => \N__26034\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_10\
        );

    \I__3408\ : InMux
    port map (
            O => \N__26031\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_11\
        );

    \I__3407\ : InMux
    port map (
            O => \N__26028\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_12\
        );

    \I__3406\ : InMux
    port map (
            O => \N__26025\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_13\
        );

    \I__3405\ : InMux
    port map (
            O => \N__26022\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_14\
        );

    \I__3404\ : InMux
    port map (
            O => \N__26019\,
            I => \bfn_10_9_0_\
        );

    \I__3403\ : InMux
    port map (
            O => \N__26016\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_16\
        );

    \I__3402\ : InMux
    port map (
            O => \N__26013\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_17\
        );

    \I__3401\ : InMux
    port map (
            O => \N__26010\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_18\
        );

    \I__3400\ : InMux
    port map (
            O => \N__26007\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_1\
        );

    \I__3399\ : InMux
    port map (
            O => \N__26004\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_2\
        );

    \I__3398\ : InMux
    port map (
            O => \N__26001\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_3\
        );

    \I__3397\ : InMux
    port map (
            O => \N__25998\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_4\
        );

    \I__3396\ : InMux
    port map (
            O => \N__25995\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_5\
        );

    \I__3395\ : InMux
    port map (
            O => \N__25992\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_6\
        );

    \I__3394\ : InMux
    port map (
            O => \N__25989\,
            I => \bfn_10_8_0_\
        );

    \I__3393\ : InMux
    port map (
            O => \N__25986\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_8\
        );

    \I__3392\ : InMux
    port map (
            O => \N__25983\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_9\
        );

    \I__3391\ : InMux
    port map (
            O => \N__25980\,
            I => \N__25977\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__25977\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__3389\ : InMux
    port map (
            O => \N__25974\,
            I => \N__25948\
        );

    \I__3388\ : InMux
    port map (
            O => \N__25973\,
            I => \N__25948\
        );

    \I__3387\ : InMux
    port map (
            O => \N__25972\,
            I => \N__25935\
        );

    \I__3386\ : InMux
    port map (
            O => \N__25971\,
            I => \N__25935\
        );

    \I__3385\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25935\
        );

    \I__3384\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25935\
        );

    \I__3383\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25922\
        );

    \I__3382\ : InMux
    port map (
            O => \N__25967\,
            I => \N__25922\
        );

    \I__3381\ : InMux
    port map (
            O => \N__25966\,
            I => \N__25922\
        );

    \I__3380\ : InMux
    port map (
            O => \N__25965\,
            I => \N__25922\
        );

    \I__3379\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25913\
        );

    \I__3378\ : InMux
    port map (
            O => \N__25963\,
            I => \N__25913\
        );

    \I__3377\ : InMux
    port map (
            O => \N__25962\,
            I => \N__25913\
        );

    \I__3376\ : InMux
    port map (
            O => \N__25961\,
            I => \N__25913\
        );

    \I__3375\ : InMux
    port map (
            O => \N__25960\,
            I => \N__25904\
        );

    \I__3374\ : InMux
    port map (
            O => \N__25959\,
            I => \N__25904\
        );

    \I__3373\ : InMux
    port map (
            O => \N__25958\,
            I => \N__25904\
        );

    \I__3372\ : InMux
    port map (
            O => \N__25957\,
            I => \N__25904\
        );

    \I__3371\ : InMux
    port map (
            O => \N__25956\,
            I => \N__25895\
        );

    \I__3370\ : InMux
    port map (
            O => \N__25955\,
            I => \N__25895\
        );

    \I__3369\ : InMux
    port map (
            O => \N__25954\,
            I => \N__25895\
        );

    \I__3368\ : InMux
    port map (
            O => \N__25953\,
            I => \N__25895\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__25948\,
            I => \N__25892\
        );

    \I__3366\ : InMux
    port map (
            O => \N__25947\,
            I => \N__25883\
        );

    \I__3365\ : InMux
    port map (
            O => \N__25946\,
            I => \N__25883\
        );

    \I__3364\ : InMux
    port map (
            O => \N__25945\,
            I => \N__25883\
        );

    \I__3363\ : InMux
    port map (
            O => \N__25944\,
            I => \N__25883\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__25935\,
            I => \N__25880\
        );

    \I__3361\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25871\
        );

    \I__3360\ : InMux
    port map (
            O => \N__25933\,
            I => \N__25871\
        );

    \I__3359\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25871\
        );

    \I__3358\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25871\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__25922\,
            I => \N__25862\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__25913\,
            I => \N__25862\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__25904\,
            I => \N__25862\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__25895\,
            I => \N__25862\
        );

    \I__3353\ : Span4Mux_v
    port map (
            O => \N__25892\,
            I => \N__25857\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__25883\,
            I => \N__25857\
        );

    \I__3351\ : Span4Mux_v
    port map (
            O => \N__25880\,
            I => \N__25848\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__25871\,
            I => \N__25848\
        );

    \I__3349\ : Span4Mux_v
    port map (
            O => \N__25862\,
            I => \N__25848\
        );

    \I__3348\ : Span4Mux_h
    port map (
            O => \N__25857\,
            I => \N__25848\
        );

    \I__3347\ : Odrv4
    port map (
            O => \N__25848\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__3346\ : InMux
    port map (
            O => \N__25845\,
            I => \N__25842\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__25842\,
            I => \N__25837\
        );

    \I__3344\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25832\
        );

    \I__3343\ : InMux
    port map (
            O => \N__25840\,
            I => \N__25832\
        );

    \I__3342\ : Span12Mux_s11_v
    port map (
            O => \N__25837\,
            I => \N__25828\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__25832\,
            I => \N__25825\
        );

    \I__3340\ : InMux
    port map (
            O => \N__25831\,
            I => \N__25822\
        );

    \I__3339\ : Span12Mux_v
    port map (
            O => \N__25828\,
            I => \N__25819\
        );

    \I__3338\ : Odrv4
    port map (
            O => \N__25825\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__25822\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__3336\ : Odrv12
    port map (
            O => \N__25819\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__3335\ : IoInMux
    port map (
            O => \N__25812\,
            I => \N__25809\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__25809\,
            I => \N__25806\
        );

    \I__3333\ : Odrv12
    port map (
            O => \N__25806\,
            I => s3_phy_c
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__25803\,
            I => \N__25798\
        );

    \I__3331\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25790\
        );

    \I__3330\ : InMux
    port map (
            O => \N__25801\,
            I => \N__25790\
        );

    \I__3329\ : InMux
    port map (
            O => \N__25798\,
            I => \N__25790\
        );

    \I__3328\ : InMux
    port map (
            O => \N__25797\,
            I => \N__25787\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__25790\,
            I => \N__25782\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__25787\,
            I => \N__25782\
        );

    \I__3325\ : Odrv4
    port map (
            O => \N__25782\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__3324\ : InMux
    port map (
            O => \N__25779\,
            I => \N__25776\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__25776\,
            I => \phase_controller_inst2.start_timer_tr_0_sqmuxa\
        );

    \I__3322\ : InMux
    port map (
            O => \N__25773\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_0\
        );

    \I__3321\ : InMux
    port map (
            O => \N__25770\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__3320\ : InMux
    port map (
            O => \N__25767\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__3319\ : InMux
    port map (
            O => \N__25764\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__3318\ : InMux
    port map (
            O => \N__25761\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__3317\ : InMux
    port map (
            O => \N__25758\,
            I => \bfn_9_22_0_\
        );

    \I__3316\ : InMux
    port map (
            O => \N__25755\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__3315\ : InMux
    port map (
            O => \N__25752\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__3314\ : InMux
    port map (
            O => \N__25749\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__3313\ : InMux
    port map (
            O => \N__25746\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__3312\ : InMux
    port map (
            O => \N__25743\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__3311\ : InMux
    port map (
            O => \N__25740\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__3310\ : InMux
    port map (
            O => \N__25737\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__3309\ : InMux
    port map (
            O => \N__25734\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__3308\ : InMux
    port map (
            O => \N__25731\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__3307\ : InMux
    port map (
            O => \N__25728\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__3306\ : InMux
    port map (
            O => \N__25725\,
            I => \bfn_9_21_0_\
        );

    \I__3305\ : InMux
    port map (
            O => \N__25722\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__3304\ : InMux
    port map (
            O => \N__25719\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__3303\ : InMux
    port map (
            O => \N__25716\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__3302\ : InMux
    port map (
            O => \N__25713\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__3301\ : InMux
    port map (
            O => \N__25710\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__3300\ : InMux
    port map (
            O => \N__25707\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__3299\ : InMux
    port map (
            O => \N__25704\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__3298\ : InMux
    port map (
            O => \N__25701\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__3297\ : InMux
    port map (
            O => \N__25698\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__3296\ : InMux
    port map (
            O => \N__25695\,
            I => \bfn_9_20_0_\
        );

    \I__3295\ : InMux
    port map (
            O => \N__25692\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__3294\ : InMux
    port map (
            O => \N__25689\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__3293\ : InMux
    port map (
            O => \N__25686\,
            I => \N__25683\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__25683\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__3291\ : CascadeMux
    port map (
            O => \N__25680\,
            I => \N__25677\
        );

    \I__3290\ : InMux
    port map (
            O => \N__25677\,
            I => \N__25674\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__25674\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__25671\,
            I => \N__25668\
        );

    \I__3287\ : InMux
    port map (
            O => \N__25668\,
            I => \N__25665\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__25665\,
            I => \N__25662\
        );

    \I__3285\ : Span4Mux_v
    port map (
            O => \N__25662\,
            I => \N__25658\
        );

    \I__3284\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25653\
        );

    \I__3283\ : Span4Mux_v
    port map (
            O => \N__25658\,
            I => \N__25650\
        );

    \I__3282\ : InMux
    port map (
            O => \N__25657\,
            I => \N__25647\
        );

    \I__3281\ : InMux
    port map (
            O => \N__25656\,
            I => \N__25644\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__25653\,
            I => \N__25641\
        );

    \I__3279\ : Odrv4
    port map (
            O => \N__25650\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__25647\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__25644\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__3276\ : Odrv12
    port map (
            O => \N__25641\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__25632\,
            I => \N__25629\
        );

    \I__3274\ : InMux
    port map (
            O => \N__25629\,
            I => \N__25626\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__25626\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__3272\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25620\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__25620\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\
        );

    \I__3270\ : CascadeMux
    port map (
            O => \N__25617\,
            I => \N__25614\
        );

    \I__3269\ : InMux
    port map (
            O => \N__25614\,
            I => \N__25611\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__25611\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__3267\ : InMux
    port map (
            O => \N__25608\,
            I => \N__25605\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__25605\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__3265\ : CascadeMux
    port map (
            O => \N__25602\,
            I => \N__25599\
        );

    \I__3264\ : InMux
    port map (
            O => \N__25599\,
            I => \N__25596\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__25596\,
            I => \N__25593\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__25593\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\
        );

    \I__3261\ : InMux
    port map (
            O => \N__25590\,
            I => \bfn_9_19_0_\
        );

    \I__3260\ : InMux
    port map (
            O => \N__25587\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__25584\,
            I => \N__25581\
        );

    \I__3258\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25578\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__25578\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__3256\ : InMux
    port map (
            O => \N__25575\,
            I => \N__25572\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__25572\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__3254\ : InMux
    port map (
            O => \N__25569\,
            I => \N__25566\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__25566\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__3252\ : InMux
    port map (
            O => \N__25563\,
            I => \N__25560\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__25560\,
            I => \N__25557\
        );

    \I__3250\ : Span4Mux_h
    port map (
            O => \N__25557\,
            I => \N__25554\
        );

    \I__3249\ : Odrv4
    port map (
            O => \N__25554\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__3248\ : InMux
    port map (
            O => \N__25551\,
            I => \N__25548\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__25548\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__25545\,
            I => \N__25542\
        );

    \I__3245\ : InMux
    port map (
            O => \N__25542\,
            I => \N__25539\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__25539\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__25536\,
            I => \N__25533\
        );

    \I__3242\ : InMux
    port map (
            O => \N__25533\,
            I => \N__25530\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__25530\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__3240\ : CascadeMux
    port map (
            O => \N__25527\,
            I => \N__25524\
        );

    \I__3239\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25521\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__25521\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__3237\ : CascadeMux
    port map (
            O => \N__25518\,
            I => \N__25515\
        );

    \I__3236\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25512\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__25512\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\
        );

    \I__3234\ : InMux
    port map (
            O => \N__25509\,
            I => \N__25506\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__25506\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__3232\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25500\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__25500\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__3230\ : InMux
    port map (
            O => \N__25497\,
            I => \N__25494\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__25494\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__3228\ : InMux
    port map (
            O => \N__25491\,
            I => \N__25488\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__25488\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__3226\ : InMux
    port map (
            O => \N__25485\,
            I => \N__25482\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__25482\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__25479\,
            I => \N__25476\
        );

    \I__3223\ : InMux
    port map (
            O => \N__25476\,
            I => \N__25473\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__25473\,
            I => \N__25470\
        );

    \I__3221\ : Span4Mux_v
    port map (
            O => \N__25470\,
            I => \N__25467\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__25467\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\
        );

    \I__3219\ : InMux
    port map (
            O => \N__25464\,
            I => \N__25461\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__25461\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__25458\,
            I => \N__25455\
        );

    \I__3216\ : InMux
    port map (
            O => \N__25455\,
            I => \N__25452\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__25452\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__3214\ : InMux
    port map (
            O => \N__25449\,
            I => \N__25446\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__25446\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__3212\ : CascadeMux
    port map (
            O => \N__25443\,
            I => \N__25440\
        );

    \I__3211\ : InMux
    port map (
            O => \N__25440\,
            I => \N__25437\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__25437\,
            I => \N__25434\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__25434\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\
        );

    \I__3208\ : InMux
    port map (
            O => \N__25431\,
            I => \N__25428\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__25428\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__25425\,
            I => \N__25422\
        );

    \I__3205\ : InMux
    port map (
            O => \N__25422\,
            I => \N__25419\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__25419\,
            I => \N__25416\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__25416\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__25413\,
            I => \N__25410\
        );

    \I__3201\ : InMux
    port map (
            O => \N__25410\,
            I => \N__25407\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__25407\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__3199\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25401\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__25401\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__3197\ : InMux
    port map (
            O => \N__25398\,
            I => \N__25395\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__25395\,
            I => \N__25392\
        );

    \I__3195\ : Span4Mux_v
    port map (
            O => \N__25392\,
            I => \N__25389\
        );

    \I__3194\ : Odrv4
    port map (
            O => \N__25389\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__25386\,
            I => \N__25383\
        );

    \I__3192\ : InMux
    port map (
            O => \N__25383\,
            I => \N__25380\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__25380\,
            I => \N__25377\
        );

    \I__3190\ : Span4Mux_h
    port map (
            O => \N__25377\,
            I => \N__25374\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__25374\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__25371\,
            I => \N__25368\
        );

    \I__3187\ : InMux
    port map (
            O => \N__25368\,
            I => \N__25365\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__25365\,
            I => \N__25362\
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__25362\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__25359\,
            I => \N__25356\
        );

    \I__3183\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25353\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__25353\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__3181\ : InMux
    port map (
            O => \N__25350\,
            I => \N__25347\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__25347\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__25344\,
            I => \N__25341\
        );

    \I__3178\ : InMux
    port map (
            O => \N__25341\,
            I => \N__25338\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__25338\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__3176\ : InMux
    port map (
            O => \N__25335\,
            I => \N__25332\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__25332\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\
        );

    \I__3174\ : InMux
    port map (
            O => \N__25329\,
            I => \N__25326\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__25326\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__25323\,
            I => \N__25320\
        );

    \I__3171\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25317\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__25317\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\
        );

    \I__3169\ : InMux
    port map (
            O => \N__25314\,
            I => \N__25311\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__25311\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\
        );

    \I__3167\ : CascadeMux
    port map (
            O => \N__25308\,
            I => \N__25305\
        );

    \I__3166\ : InMux
    port map (
            O => \N__25305\,
            I => \N__25302\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__25302\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__25299\,
            I => \N__25296\
        );

    \I__3163\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25293\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__25293\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\
        );

    \I__3161\ : InMux
    port map (
            O => \N__25290\,
            I => \N__25287\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__25287\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__3159\ : InMux
    port map (
            O => \N__25284\,
            I => \N__25281\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__25281\,
            I => \N__25277\
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__25280\,
            I => \N__25274\
        );

    \I__3156\ : Span12Mux_s8_v
    port map (
            O => \N__25277\,
            I => \N__25269\
        );

    \I__3155\ : InMux
    port map (
            O => \N__25274\,
            I => \N__25266\
        );

    \I__3154\ : InMux
    port map (
            O => \N__25273\,
            I => \N__25263\
        );

    \I__3153\ : InMux
    port map (
            O => \N__25272\,
            I => \N__25260\
        );

    \I__3152\ : Span12Mux_v
    port map (
            O => \N__25269\,
            I => \N__25257\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__25266\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__25263\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__25260\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3148\ : Odrv12
    port map (
            O => \N__25257\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3147\ : InMux
    port map (
            O => \N__25248\,
            I => \N__25245\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__25245\,
            I => \N__25242\
        );

    \I__3145\ : Span4Mux_v
    port map (
            O => \N__25242\,
            I => \N__25237\
        );

    \I__3144\ : InMux
    port map (
            O => \N__25241\,
            I => \N__25234\
        );

    \I__3143\ : InMux
    port map (
            O => \N__25240\,
            I => \N__25231\
        );

    \I__3142\ : Sp12to4
    port map (
            O => \N__25237\,
            I => \N__25224\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__25234\,
            I => \N__25224\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__25231\,
            I => \N__25224\
        );

    \I__3139\ : Span12Mux_h
    port map (
            O => \N__25224\,
            I => \N__25221\
        );

    \I__3138\ : Odrv12
    port map (
            O => \N__25221\,
            I => il_min_comp2_c
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__25218\,
            I => \N__25213\
        );

    \I__3136\ : InMux
    port map (
            O => \N__25217\,
            I => \N__25208\
        );

    \I__3135\ : InMux
    port map (
            O => \N__25216\,
            I => \N__25208\
        );

    \I__3134\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25205\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__25208\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__25205\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__25200\,
            I => \N__25197\
        );

    \I__3130\ : InMux
    port map (
            O => \N__25197\,
            I => \N__25193\
        );

    \I__3129\ : InMux
    port map (
            O => \N__25196\,
            I => \N__25190\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__25193\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__25190\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__25185\,
            I => \N__25182\
        );

    \I__3125\ : InMux
    port map (
            O => \N__25182\,
            I => \N__25179\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__25179\,
            I => \phase_controller_inst2.stoper_tr.un4_start_0\
        );

    \I__3123\ : InMux
    port map (
            O => \N__25176\,
            I => \N__25173\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__25173\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\
        );

    \I__3121\ : InMux
    port map (
            O => \N__25170\,
            I => \N__25167\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__25167\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__25164\,
            I => \N__25161\
        );

    \I__3118\ : InMux
    port map (
            O => \N__25161\,
            I => \N__25158\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__25158\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__3116\ : InMux
    port map (
            O => \N__25155\,
            I => \N__25152\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__25152\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\
        );

    \I__3114\ : InMux
    port map (
            O => \N__25149\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__3113\ : InMux
    port map (
            O => \N__25146\,
            I => \N__25143\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__25143\,
            I => \N__25140\
        );

    \I__3111\ : Span4Mux_h
    port map (
            O => \N__25140\,
            I => \N__25137\
        );

    \I__3110\ : Span4Mux_v
    port map (
            O => \N__25137\,
            I => \N__25134\
        );

    \I__3109\ : Odrv4
    port map (
            O => \N__25134\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__3108\ : InMux
    port map (
            O => \N__25131\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__3107\ : CascadeMux
    port map (
            O => \N__25128\,
            I => \N__25125\
        );

    \I__3106\ : InMux
    port map (
            O => \N__25125\,
            I => \N__25122\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__25122\,
            I => \N__25119\
        );

    \I__3104\ : Span4Mux_v
    port map (
            O => \N__25119\,
            I => \N__25116\
        );

    \I__3103\ : Odrv4
    port map (
            O => \N__25116\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__3102\ : InMux
    port map (
            O => \N__25113\,
            I => \N__25110\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__25110\,
            I => \N__25107\
        );

    \I__3100\ : Span12Mux_v
    port map (
            O => \N__25107\,
            I => \N__25104\
        );

    \I__3099\ : Odrv12
    port map (
            O => \N__25104\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__3098\ : InMux
    port map (
            O => \N__25101\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__3097\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25095\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__25095\,
            I => \N__25092\
        );

    \I__3095\ : Span4Mux_h
    port map (
            O => \N__25092\,
            I => \N__25089\
        );

    \I__3094\ : Sp12to4
    port map (
            O => \N__25089\,
            I => \N__25086\
        );

    \I__3093\ : Odrv12
    port map (
            O => \N__25086\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__3092\ : InMux
    port map (
            O => \N__25083\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__3091\ : InMux
    port map (
            O => \N__25080\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__3090\ : InMux
    port map (
            O => \N__25077\,
            I => \N__25074\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__25074\,
            I => \N__25071\
        );

    \I__3088\ : Span12Mux_v
    port map (
            O => \N__25071\,
            I => \N__25068\
        );

    \I__3087\ : Odrv12
    port map (
            O => \N__25068\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__25065\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\
        );

    \I__3085\ : InMux
    port map (
            O => \N__25062\,
            I => \N__25059\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__25059\,
            I => \N__25055\
        );

    \I__3083\ : InMux
    port map (
            O => \N__25058\,
            I => \N__25052\
        );

    \I__3082\ : Span12Mux_v
    port map (
            O => \N__25055\,
            I => \N__25047\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__25052\,
            I => \N__25047\
        );

    \I__3080\ : Odrv12
    port map (
            O => \N__25047\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__3079\ : IoInMux
    port map (
            O => \N__25044\,
            I => \N__25041\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__25041\,
            I => \N__25038\
        );

    \I__3077\ : Odrv12
    port map (
            O => \N__25038\,
            I => s4_phy_c
        );

    \I__3076\ : InMux
    port map (
            O => \N__25035\,
            I => \N__25032\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__25032\,
            I => \N__25029\
        );

    \I__3074\ : Odrv4
    port map (
            O => \N__25029\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\
        );

    \I__3073\ : InMux
    port map (
            O => \N__25026\,
            I => \N__25023\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__25023\,
            I => \N__25020\
        );

    \I__3071\ : Span4Mux_h
    port map (
            O => \N__25020\,
            I => \N__25017\
        );

    \I__3070\ : Odrv4
    port map (
            O => \N__25017\,
            I => \current_shift_inst.un38_control_input_0_s1_19\
        );

    \I__3069\ : InMux
    port map (
            O => \N__25014\,
            I => \current_shift_inst.un38_control_input_cry_18_s1\
        );

    \I__3068\ : InMux
    port map (
            O => \N__25011\,
            I => \N__25008\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__25008\,
            I => \N__25005\
        );

    \I__3066\ : Sp12to4
    port map (
            O => \N__25005\,
            I => \N__25002\
        );

    \I__3065\ : Odrv12
    port map (
            O => \N__25002\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__3064\ : InMux
    port map (
            O => \N__24999\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__3063\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24993\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__24993\,
            I => \N__24990\
        );

    \I__3061\ : Span4Mux_h
    port map (
            O => \N__24990\,
            I => \N__24987\
        );

    \I__3060\ : Sp12to4
    port map (
            O => \N__24987\,
            I => \N__24984\
        );

    \I__3059\ : Odrv12
    port map (
            O => \N__24984\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__3058\ : InMux
    port map (
            O => \N__24981\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__3057\ : InMux
    port map (
            O => \N__24978\,
            I => \N__24975\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__24975\,
            I => \N__24972\
        );

    \I__3055\ : Span4Mux_v
    port map (
            O => \N__24972\,
            I => \N__24969\
        );

    \I__3054\ : Odrv4
    port map (
            O => \N__24969\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__3053\ : InMux
    port map (
            O => \N__24966\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__3052\ : InMux
    port map (
            O => \N__24963\,
            I => \N__24960\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__24960\,
            I => \N__24957\
        );

    \I__3050\ : Span4Mux_h
    port map (
            O => \N__24957\,
            I => \N__24954\
        );

    \I__3049\ : Span4Mux_v
    port map (
            O => \N__24954\,
            I => \N__24951\
        );

    \I__3048\ : Span4Mux_v
    port map (
            O => \N__24951\,
            I => \N__24948\
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__24948\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__3046\ : InMux
    port map (
            O => \N__24945\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__3045\ : InMux
    port map (
            O => \N__24942\,
            I => \N__24939\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__24939\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__3043\ : InMux
    port map (
            O => \N__24936\,
            I => \N__24933\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__24933\,
            I => \N__24930\
        );

    \I__3041\ : Span4Mux_v
    port map (
            O => \N__24930\,
            I => \N__24927\
        );

    \I__3040\ : Odrv4
    port map (
            O => \N__24927\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__3039\ : InMux
    port map (
            O => \N__24924\,
            I => \bfn_8_22_0_\
        );

    \I__3038\ : InMux
    port map (
            O => \N__24921\,
            I => \N__24918\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__24918\,
            I => \N__24915\
        );

    \I__3036\ : Span4Mux_h
    port map (
            O => \N__24915\,
            I => \N__24912\
        );

    \I__3035\ : Span4Mux_v
    port map (
            O => \N__24912\,
            I => \N__24909\
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__24909\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__3033\ : InMux
    port map (
            O => \N__24906\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__3032\ : InMux
    port map (
            O => \N__24903\,
            I => \N__24900\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__24900\,
            I => \N__24897\
        );

    \I__3030\ : Span4Mux_h
    port map (
            O => \N__24897\,
            I => \N__24894\
        );

    \I__3029\ : Span4Mux_v
    port map (
            O => \N__24894\,
            I => \N__24891\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__24891\,
            I => \N__24888\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__24888\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__3026\ : InMux
    port map (
            O => \N__24885\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__3025\ : InMux
    port map (
            O => \N__24882\,
            I => \N__24879\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__24879\,
            I => \N__24876\
        );

    \I__3023\ : Span4Mux_h
    port map (
            O => \N__24876\,
            I => \N__24873\
        );

    \I__3022\ : Span4Mux_v
    port map (
            O => \N__24873\,
            I => \N__24870\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__24870\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__24867\,
            I => \N__24864\
        );

    \I__3019\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24861\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__24861\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\
        );

    \I__3017\ : InMux
    port map (
            O => \N__24858\,
            I => \N__24855\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__24855\,
            I => \N__24852\
        );

    \I__3015\ : Span4Mux_h
    port map (
            O => \N__24852\,
            I => \N__24849\
        );

    \I__3014\ : Span4Mux_v
    port map (
            O => \N__24849\,
            I => \N__24846\
        );

    \I__3013\ : Odrv4
    port map (
            O => \N__24846\,
            I => \current_shift_inst.un38_control_input_0_s1_11\
        );

    \I__3012\ : InMux
    port map (
            O => \N__24843\,
            I => \current_shift_inst.un38_control_input_cry_10_s1\
        );

    \I__3011\ : InMux
    port map (
            O => \N__24840\,
            I => \N__24837\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__24837\,
            I => \N__24834\
        );

    \I__3009\ : Sp12to4
    port map (
            O => \N__24834\,
            I => \N__24831\
        );

    \I__3008\ : Odrv12
    port map (
            O => \N__24831\,
            I => \current_shift_inst.un38_control_input_0_s1_12\
        );

    \I__3007\ : InMux
    port map (
            O => \N__24828\,
            I => \current_shift_inst.un38_control_input_cry_11_s1\
        );

    \I__3006\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24822\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__24822\,
            I => \N__24819\
        );

    \I__3004\ : Span12Mux_s8_h
    port map (
            O => \N__24819\,
            I => \N__24816\
        );

    \I__3003\ : Odrv12
    port map (
            O => \N__24816\,
            I => \current_shift_inst.un38_control_input_0_s1_13\
        );

    \I__3002\ : InMux
    port map (
            O => \N__24813\,
            I => \current_shift_inst.un38_control_input_cry_12_s1\
        );

    \I__3001\ : InMux
    port map (
            O => \N__24810\,
            I => \N__24807\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__24807\,
            I => \N__24804\
        );

    \I__2999\ : Span4Mux_v
    port map (
            O => \N__24804\,
            I => \N__24801\
        );

    \I__2998\ : Span4Mux_v
    port map (
            O => \N__24801\,
            I => \N__24798\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__24798\,
            I => \current_shift_inst.un38_control_input_0_s1_14\
        );

    \I__2996\ : InMux
    port map (
            O => \N__24795\,
            I => \current_shift_inst.un38_control_input_cry_13_s1\
        );

    \I__2995\ : InMux
    port map (
            O => \N__24792\,
            I => \N__24789\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__24789\,
            I => \N__24786\
        );

    \I__2993\ : Sp12to4
    port map (
            O => \N__24786\,
            I => \N__24783\
        );

    \I__2992\ : Span12Mux_v
    port map (
            O => \N__24783\,
            I => \N__24780\
        );

    \I__2991\ : Odrv12
    port map (
            O => \N__24780\,
            I => \current_shift_inst.un38_control_input_0_s1_15\
        );

    \I__2990\ : InMux
    port map (
            O => \N__24777\,
            I => \current_shift_inst.un38_control_input_cry_14_s1\
        );

    \I__2989\ : InMux
    port map (
            O => \N__24774\,
            I => \N__24771\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__24771\,
            I => \N__24768\
        );

    \I__2987\ : Span12Mux_v
    port map (
            O => \N__24768\,
            I => \N__24765\
        );

    \I__2986\ : Odrv12
    port map (
            O => \N__24765\,
            I => \current_shift_inst.un38_control_input_0_s1_16\
        );

    \I__2985\ : InMux
    port map (
            O => \N__24762\,
            I => \bfn_8_21_0_\
        );

    \I__2984\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24756\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__24756\,
            I => \N__24753\
        );

    \I__2982\ : Span4Mux_v
    port map (
            O => \N__24753\,
            I => \N__24750\
        );

    \I__2981\ : Span4Mux_v
    port map (
            O => \N__24750\,
            I => \N__24747\
        );

    \I__2980\ : Odrv4
    port map (
            O => \N__24747\,
            I => \current_shift_inst.un38_control_input_0_s1_17\
        );

    \I__2979\ : InMux
    port map (
            O => \N__24744\,
            I => \current_shift_inst.un38_control_input_cry_16_s1\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__24741\,
            I => \N__24738\
        );

    \I__2977\ : InMux
    port map (
            O => \N__24738\,
            I => \N__24735\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__24735\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\
        );

    \I__2975\ : InMux
    port map (
            O => \N__24732\,
            I => \N__24729\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__24729\,
            I => \N__24726\
        );

    \I__2973\ : Span4Mux_v
    port map (
            O => \N__24726\,
            I => \N__24723\
        );

    \I__2972\ : Odrv4
    port map (
            O => \N__24723\,
            I => \current_shift_inst.un38_control_input_0_s1_18\
        );

    \I__2971\ : InMux
    port map (
            O => \N__24720\,
            I => \current_shift_inst.un38_control_input_cry_17_s1\
        );

    \I__2970\ : InMux
    port map (
            O => \N__24717\,
            I => \N__24714\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__24714\,
            I => \N__24711\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__24711\,
            I => \current_shift_inst.un38_control_input_0_s1_3\
        );

    \I__2967\ : InMux
    port map (
            O => \N__24708\,
            I => \current_shift_inst.un38_control_input_cry_2_s1\
        );

    \I__2966\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24702\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__24702\,
            I => \N__24699\
        );

    \I__2964\ : Odrv4
    port map (
            O => \N__24699\,
            I => \current_shift_inst.un38_control_input_0_s1_4\
        );

    \I__2963\ : InMux
    port map (
            O => \N__24696\,
            I => \current_shift_inst.un38_control_input_cry_3_s1\
        );

    \I__2962\ : InMux
    port map (
            O => \N__24693\,
            I => \N__24690\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__24690\,
            I => \N__24687\
        );

    \I__2960\ : Span12Mux_s8_h
    port map (
            O => \N__24687\,
            I => \N__24684\
        );

    \I__2959\ : Odrv12
    port map (
            O => \N__24684\,
            I => \current_shift_inst.un38_control_input_0_s1_5\
        );

    \I__2958\ : InMux
    port map (
            O => \N__24681\,
            I => \current_shift_inst.un38_control_input_cry_4_s1\
        );

    \I__2957\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24675\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__24675\,
            I => \N__24672\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__24672\,
            I => \current_shift_inst.un38_control_input_0_s1_6\
        );

    \I__2954\ : InMux
    port map (
            O => \N__24669\,
            I => \current_shift_inst.un38_control_input_cry_5_s1\
        );

    \I__2953\ : InMux
    port map (
            O => \N__24666\,
            I => \N__24663\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__24663\,
            I => \N__24660\
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__24660\,
            I => \current_shift_inst.un38_control_input_0_s1_7\
        );

    \I__2950\ : InMux
    port map (
            O => \N__24657\,
            I => \current_shift_inst.un38_control_input_cry_6_s1\
        );

    \I__2949\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24651\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__24651\,
            I => \N__24648\
        );

    \I__2947\ : Span12Mux_v
    port map (
            O => \N__24648\,
            I => \N__24645\
        );

    \I__2946\ : Odrv12
    port map (
            O => \N__24645\,
            I => \current_shift_inst.un38_control_input_0_s1_8\
        );

    \I__2945\ : InMux
    port map (
            O => \N__24642\,
            I => \bfn_8_20_0_\
        );

    \I__2944\ : InMux
    port map (
            O => \N__24639\,
            I => \N__24636\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__24636\,
            I => \N__24633\
        );

    \I__2942\ : Span4Mux_h
    port map (
            O => \N__24633\,
            I => \N__24630\
        );

    \I__2941\ : Span4Mux_v
    port map (
            O => \N__24630\,
            I => \N__24627\
        );

    \I__2940\ : Odrv4
    port map (
            O => \N__24627\,
            I => \current_shift_inst.un38_control_input_0_s1_9\
        );

    \I__2939\ : InMux
    port map (
            O => \N__24624\,
            I => \current_shift_inst.un38_control_input_cry_8_s1\
        );

    \I__2938\ : InMux
    port map (
            O => \N__24621\,
            I => \N__24618\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__24618\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\
        );

    \I__2936\ : InMux
    port map (
            O => \N__24615\,
            I => \N__24612\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__24612\,
            I => \N__24609\
        );

    \I__2934\ : Span4Mux_h
    port map (
            O => \N__24609\,
            I => \N__24606\
        );

    \I__2933\ : Span4Mux_v
    port map (
            O => \N__24606\,
            I => \N__24603\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__24603\,
            I => \current_shift_inst.un38_control_input_0_s1_10\
        );

    \I__2931\ : InMux
    port map (
            O => \N__24600\,
            I => \current_shift_inst.un38_control_input_cry_9_s1\
        );

    \I__2930\ : InMux
    port map (
            O => \N__24597\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__2929\ : CascadeMux
    port map (
            O => \N__24594\,
            I => \N__24589\
        );

    \I__2928\ : InMux
    port map (
            O => \N__24593\,
            I => \N__24574\
        );

    \I__2927\ : InMux
    port map (
            O => \N__24592\,
            I => \N__24574\
        );

    \I__2926\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24569\
        );

    \I__2925\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24569\
        );

    \I__2924\ : CascadeMux
    port map (
            O => \N__24587\,
            I => \N__24566\
        );

    \I__2923\ : InMux
    port map (
            O => \N__24586\,
            I => \N__24555\
        );

    \I__2922\ : InMux
    port map (
            O => \N__24585\,
            I => \N__24544\
        );

    \I__2921\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24544\
        );

    \I__2920\ : InMux
    port map (
            O => \N__24583\,
            I => \N__24544\
        );

    \I__2919\ : InMux
    port map (
            O => \N__24582\,
            I => \N__24544\
        );

    \I__2918\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24544\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__24580\,
            I => \N__24541\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__24579\,
            I => \N__24537\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__24574\,
            I => \N__24528\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__24569\,
            I => \N__24528\
        );

    \I__2913\ : InMux
    port map (
            O => \N__24566\,
            I => \N__24515\
        );

    \I__2912\ : InMux
    port map (
            O => \N__24565\,
            I => \N__24515\
        );

    \I__2911\ : InMux
    port map (
            O => \N__24564\,
            I => \N__24515\
        );

    \I__2910\ : InMux
    port map (
            O => \N__24563\,
            I => \N__24515\
        );

    \I__2909\ : InMux
    port map (
            O => \N__24562\,
            I => \N__24515\
        );

    \I__2908\ : InMux
    port map (
            O => \N__24561\,
            I => \N__24515\
        );

    \I__2907\ : InMux
    port map (
            O => \N__24560\,
            I => \N__24512\
        );

    \I__2906\ : InMux
    port map (
            O => \N__24559\,
            I => \N__24509\
        );

    \I__2905\ : InMux
    port map (
            O => \N__24558\,
            I => \N__24506\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__24555\,
            I => \N__24501\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__24544\,
            I => \N__24501\
        );

    \I__2902\ : InMux
    port map (
            O => \N__24541\,
            I => \N__24496\
        );

    \I__2901\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24496\
        );

    \I__2900\ : InMux
    port map (
            O => \N__24537\,
            I => \N__24493\
        );

    \I__2899\ : InMux
    port map (
            O => \N__24536\,
            I => \N__24490\
        );

    \I__2898\ : InMux
    port map (
            O => \N__24535\,
            I => \N__24483\
        );

    \I__2897\ : InMux
    port map (
            O => \N__24534\,
            I => \N__24483\
        );

    \I__2896\ : InMux
    port map (
            O => \N__24533\,
            I => \N__24483\
        );

    \I__2895\ : Span4Mux_h
    port map (
            O => \N__24528\,
            I => \N__24476\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__24515\,
            I => \N__24476\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__24512\,
            I => \N__24476\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__24509\,
            I => \N__24466\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__24506\,
            I => \N__24466\
        );

    \I__2890\ : Span4Mux_v
    port map (
            O => \N__24501\,
            I => \N__24466\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__24496\,
            I => \N__24466\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__24493\,
            I => \N__24459\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__24490\,
            I => \N__24459\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__24483\,
            I => \N__24459\
        );

    \I__2885\ : Sp12to4
    port map (
            O => \N__24476\,
            I => \N__24451\
        );

    \I__2884\ : InMux
    port map (
            O => \N__24475\,
            I => \N__24448\
        );

    \I__2883\ : Span4Mux_h
    port map (
            O => \N__24466\,
            I => \N__24443\
        );

    \I__2882\ : Span4Mux_v
    port map (
            O => \N__24459\,
            I => \N__24443\
        );

    \I__2881\ : InMux
    port map (
            O => \N__24458\,
            I => \N__24432\
        );

    \I__2880\ : InMux
    port map (
            O => \N__24457\,
            I => \N__24432\
        );

    \I__2879\ : InMux
    port map (
            O => \N__24456\,
            I => \N__24432\
        );

    \I__2878\ : InMux
    port map (
            O => \N__24455\,
            I => \N__24432\
        );

    \I__2877\ : InMux
    port map (
            O => \N__24454\,
            I => \N__24432\
        );

    \I__2876\ : Span12Mux_v
    port map (
            O => \N__24451\,
            I => \N__24429\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__24448\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__24443\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__24432\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__2872\ : Odrv12
    port map (
            O => \N__24429\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__2871\ : InMux
    port map (
            O => \N__24420\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__2870\ : InMux
    port map (
            O => \N__24417\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__2869\ : InMux
    port map (
            O => \N__24414\,
            I => \N__24411\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__24411\,
            I => \N__24408\
        );

    \I__2867\ : Odrv12
    port map (
            O => \N__24408\,
            I => \current_shift_inst.control_input_axb_28\
        );

    \I__2866\ : CascadeMux
    port map (
            O => \N__24405\,
            I => \N__24402\
        );

    \I__2865\ : InMux
    port map (
            O => \N__24402\,
            I => \N__24399\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__24399\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__2863\ : InMux
    port map (
            O => \N__24396\,
            I => \N__24393\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__24393\,
            I => \N__24390\
        );

    \I__2861\ : Span4Mux_v
    port map (
            O => \N__24390\,
            I => \N__24387\
        );

    \I__2860\ : Odrv4
    port map (
            O => \N__24387\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__2859\ : InMux
    port map (
            O => \N__24384\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__2858\ : InMux
    port map (
            O => \N__24381\,
            I => \N__24378\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__24378\,
            I => \N__24375\
        );

    \I__2856\ : Odrv12
    port map (
            O => \N__24375\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__2855\ : InMux
    port map (
            O => \N__24372\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__2854\ : CascadeMux
    port map (
            O => \N__24369\,
            I => \N__24366\
        );

    \I__2853\ : InMux
    port map (
            O => \N__24366\,
            I => \N__24363\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__24363\,
            I => \N__24360\
        );

    \I__2851\ : Odrv4
    port map (
            O => \N__24360\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__2850\ : InMux
    port map (
            O => \N__24357\,
            I => \N__24354\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__24354\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__2848\ : InMux
    port map (
            O => \N__24351\,
            I => \bfn_8_14_0_\
        );

    \I__2847\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24345\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__24345\,
            I => \N__24342\
        );

    \I__2845\ : Odrv12
    port map (
            O => \N__24342\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__2844\ : InMux
    port map (
            O => \N__24339\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__2843\ : InMux
    port map (
            O => \N__24336\,
            I => \N__24333\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__24333\,
            I => \N__24330\
        );

    \I__2841\ : Odrv12
    port map (
            O => \N__24330\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__2840\ : InMux
    port map (
            O => \N__24327\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__2839\ : InMux
    port map (
            O => \N__24324\,
            I => \N__24321\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__24321\,
            I => \N__24318\
        );

    \I__2837\ : Span4Mux_h
    port map (
            O => \N__24318\,
            I => \N__24315\
        );

    \I__2836\ : Odrv4
    port map (
            O => \N__24315\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__2835\ : InMux
    port map (
            O => \N__24312\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__2834\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24306\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__24306\,
            I => \N__24303\
        );

    \I__2832\ : Odrv12
    port map (
            O => \N__24303\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__2831\ : InMux
    port map (
            O => \N__24300\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__2830\ : InMux
    port map (
            O => \N__24297\,
            I => \N__24294\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__24294\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__2828\ : InMux
    port map (
            O => \N__24291\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__2827\ : InMux
    port map (
            O => \N__24288\,
            I => \N__24285\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__24285\,
            I => \N__24282\
        );

    \I__2825\ : Span4Mux_h
    port map (
            O => \N__24282\,
            I => \N__24279\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__24279\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__2823\ : InMux
    port map (
            O => \N__24276\,
            I => \N__24273\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__24273\,
            I => \current_shift_inst.un38_control_input_0_s0_14\
        );

    \I__2821\ : InMux
    port map (
            O => \N__24270\,
            I => \current_shift_inst.un38_control_input_cry_13_s0\
        );

    \I__2820\ : InMux
    port map (
            O => \N__24267\,
            I => \N__24264\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__24264\,
            I => \N__24261\
        );

    \I__2818\ : Span4Mux_h
    port map (
            O => \N__24261\,
            I => \N__24258\
        );

    \I__2817\ : Odrv4
    port map (
            O => \N__24258\,
            I => \current_shift_inst.un38_control_input_0_s0_15\
        );

    \I__2816\ : InMux
    port map (
            O => \N__24255\,
            I => \current_shift_inst.un38_control_input_cry_14_s0\
        );

    \I__2815\ : InMux
    port map (
            O => \N__24252\,
            I => \N__24249\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__24249\,
            I => \N__24246\
        );

    \I__2813\ : Odrv12
    port map (
            O => \N__24246\,
            I => \current_shift_inst.un38_control_input_0_s0_16\
        );

    \I__2812\ : InMux
    port map (
            O => \N__24243\,
            I => \bfn_8_13_0_\
        );

    \I__2811\ : InMux
    port map (
            O => \N__24240\,
            I => \N__24237\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__24237\,
            I => \current_shift_inst.un38_control_input_0_s0_17\
        );

    \I__2809\ : InMux
    port map (
            O => \N__24234\,
            I => \current_shift_inst.un38_control_input_cry_16_s0\
        );

    \I__2808\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24228\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__24228\,
            I => \N__24225\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__24225\,
            I => \current_shift_inst.un38_control_input_0_s0_18\
        );

    \I__2805\ : InMux
    port map (
            O => \N__24222\,
            I => \current_shift_inst.un38_control_input_cry_17_s0\
        );

    \I__2804\ : InMux
    port map (
            O => \N__24219\,
            I => \N__24216\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__24216\,
            I => \N__24213\
        );

    \I__2802\ : Span4Mux_v
    port map (
            O => \N__24213\,
            I => \N__24210\
        );

    \I__2801\ : Odrv4
    port map (
            O => \N__24210\,
            I => \current_shift_inst.un38_control_input_0_s0_19\
        );

    \I__2800\ : InMux
    port map (
            O => \N__24207\,
            I => \current_shift_inst.un38_control_input_cry_18_s0\
        );

    \I__2799\ : InMux
    port map (
            O => \N__24204\,
            I => \N__24201\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__24201\,
            I => \N__24198\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__24198\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__2796\ : InMux
    port map (
            O => \N__24195\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__2795\ : InMux
    port map (
            O => \N__24192\,
            I => \N__24189\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__24189\,
            I => \N__24186\
        );

    \I__2793\ : Odrv12
    port map (
            O => \N__24186\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__2792\ : InMux
    port map (
            O => \N__24183\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__2791\ : InMux
    port map (
            O => \N__24180\,
            I => \current_shift_inst.un38_control_input_cry_4_s0\
        );

    \I__2790\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24174\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__24174\,
            I => \N__24171\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__24171\,
            I => \N__24168\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__24168\,
            I => \current_shift_inst.un38_control_input_0_s0_6\
        );

    \I__2786\ : InMux
    port map (
            O => \N__24165\,
            I => \current_shift_inst.un38_control_input_cry_5_s0\
        );

    \I__2785\ : InMux
    port map (
            O => \N__24162\,
            I => \N__24159\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__24159\,
            I => \N__24156\
        );

    \I__2783\ : Span4Mux_v
    port map (
            O => \N__24156\,
            I => \N__24153\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__24153\,
            I => \current_shift_inst.un38_control_input_0_s0_7\
        );

    \I__2781\ : InMux
    port map (
            O => \N__24150\,
            I => \current_shift_inst.un38_control_input_cry_6_s0\
        );

    \I__2780\ : InMux
    port map (
            O => \N__24147\,
            I => \N__24144\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__24144\,
            I => \N__24141\
        );

    \I__2778\ : Odrv12
    port map (
            O => \N__24141\,
            I => \current_shift_inst.un38_control_input_0_s0_8\
        );

    \I__2777\ : InMux
    port map (
            O => \N__24138\,
            I => \bfn_8_12_0_\
        );

    \I__2776\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24132\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__24132\,
            I => \N__24129\
        );

    \I__2774\ : Odrv12
    port map (
            O => \N__24129\,
            I => \current_shift_inst.un38_control_input_0_s0_9\
        );

    \I__2773\ : InMux
    port map (
            O => \N__24126\,
            I => \current_shift_inst.un38_control_input_cry_8_s0\
        );

    \I__2772\ : InMux
    port map (
            O => \N__24123\,
            I => \N__24120\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__24120\,
            I => \N__24117\
        );

    \I__2770\ : Odrv12
    port map (
            O => \N__24117\,
            I => \current_shift_inst.un38_control_input_0_s0_10\
        );

    \I__2769\ : InMux
    port map (
            O => \N__24114\,
            I => \current_shift_inst.un38_control_input_cry_9_s0\
        );

    \I__2768\ : InMux
    port map (
            O => \N__24111\,
            I => \N__24108\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__24108\,
            I => \N__24105\
        );

    \I__2766\ : Odrv12
    port map (
            O => \N__24105\,
            I => \current_shift_inst.un38_control_input_0_s0_11\
        );

    \I__2765\ : InMux
    port map (
            O => \N__24102\,
            I => \current_shift_inst.un38_control_input_cry_10_s0\
        );

    \I__2764\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24096\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__24096\,
            I => \current_shift_inst.un38_control_input_0_s0_12\
        );

    \I__2762\ : InMux
    port map (
            O => \N__24093\,
            I => \current_shift_inst.un38_control_input_cry_11_s0\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__24090\,
            I => \N__24087\
        );

    \I__2760\ : InMux
    port map (
            O => \N__24087\,
            I => \N__24084\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__24084\,
            I => \N__24081\
        );

    \I__2758\ : Span4Mux_v
    port map (
            O => \N__24081\,
            I => \N__24078\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__24078\,
            I => \current_shift_inst.un38_control_input_0_s0_13\
        );

    \I__2756\ : InMux
    port map (
            O => \N__24075\,
            I => \current_shift_inst.un38_control_input_cry_12_s0\
        );

    \I__2755\ : InMux
    port map (
            O => \N__24072\,
            I => \N__24063\
        );

    \I__2754\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24063\
        );

    \I__2753\ : InMux
    port map (
            O => \N__24070\,
            I => \N__24063\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__24063\,
            I => \phase_controller_inst2.stateZ0Z_4\
        );

    \I__2751\ : CascadeMux
    port map (
            O => \N__24060\,
            I => \N__24055\
        );

    \I__2750\ : CascadeMux
    port map (
            O => \N__24059\,
            I => \N__24052\
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__24058\,
            I => \N__24049\
        );

    \I__2748\ : InMux
    port map (
            O => \N__24055\,
            I => \N__24042\
        );

    \I__2747\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24042\
        );

    \I__2746\ : InMux
    port map (
            O => \N__24049\,
            I => \N__24042\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__24042\,
            I => \phase_controller_inst2.start_flagZ0\
        );

    \I__2744\ : InMux
    port map (
            O => \N__24039\,
            I => \N__24036\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__24036\,
            I => \phase_controller_inst2.state_ns_0_0_1\
        );

    \I__2742\ : InMux
    port map (
            O => \N__24033\,
            I => \N__24030\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__24030\,
            I => \N__24027\
        );

    \I__2740\ : Span4Mux_v
    port map (
            O => \N__24027\,
            I => \N__24024\
        );

    \I__2739\ : Odrv4
    port map (
            O => \N__24024\,
            I => \current_shift_inst.un38_control_input_0_s0_3\
        );

    \I__2738\ : InMux
    port map (
            O => \N__24021\,
            I => \current_shift_inst.un38_control_input_cry_2_s0\
        );

    \I__2737\ : InMux
    port map (
            O => \N__24018\,
            I => \N__24015\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__24015\,
            I => \N__24012\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__24012\,
            I => \N__24009\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__24009\,
            I => \current_shift_inst.un38_control_input_0_s0_4\
        );

    \I__2733\ : InMux
    port map (
            O => \N__24006\,
            I => \current_shift_inst.un38_control_input_cry_3_s0\
        );

    \I__2732\ : InMux
    port map (
            O => \N__24003\,
            I => \N__24000\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__24000\,
            I => \N__23997\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__23997\,
            I => \N__23994\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__23994\,
            I => \current_shift_inst.un38_control_input_0_s0_5\
        );

    \I__2728\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23987\
        );

    \I__2727\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23984\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__23987\,
            I => \N__23981\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__23984\,
            I => \N__23978\
        );

    \I__2724\ : Span4Mux_v
    port map (
            O => \N__23981\,
            I => \N__23975\
        );

    \I__2723\ : Span4Mux_v
    port map (
            O => \N__23978\,
            I => \N__23972\
        );

    \I__2722\ : Span4Mux_v
    port map (
            O => \N__23975\,
            I => \N__23969\
        );

    \I__2721\ : Span4Mux_h
    port map (
            O => \N__23972\,
            I => \N__23966\
        );

    \I__2720\ : Odrv4
    port map (
            O => \N__23969\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__23966\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__2718\ : InMux
    port map (
            O => \N__23961\,
            I => \N__23958\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__23958\,
            I => \N__23954\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__23957\,
            I => \N__23951\
        );

    \I__2715\ : Span4Mux_v
    port map (
            O => \N__23954\,
            I => \N__23947\
        );

    \I__2714\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23942\
        );

    \I__2713\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23942\
        );

    \I__2712\ : Sp12to4
    port map (
            O => \N__23947\,
            I => \N__23937\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__23942\,
            I => \N__23937\
        );

    \I__2710\ : Span12Mux_h
    port map (
            O => \N__23937\,
            I => \N__23934\
        );

    \I__2709\ : Odrv12
    port map (
            O => \N__23934\,
            I => il_max_comp2_c
        );

    \I__2708\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23928\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__23928\,
            I => \N__23925\
        );

    \I__2706\ : Span4Mux_h
    port map (
            O => \N__23925\,
            I => \N__23922\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__23922\,
            I => \N__23919\
        );

    \I__2704\ : Odrv4
    port map (
            O => \N__23919\,
            I => \current_shift_inst.control_input_axb_19\
        );

    \I__2703\ : InMux
    port map (
            O => \N__23916\,
            I => \N__23912\
        );

    \I__2702\ : InMux
    port map (
            O => \N__23915\,
            I => \N__23909\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__23912\,
            I => \N__23906\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__23909\,
            I => \N__23903\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__23906\,
            I => \N__23900\
        );

    \I__2698\ : Span4Mux_s1_h
    port map (
            O => \N__23903\,
            I => \N__23897\
        );

    \I__2697\ : Span4Mux_v
    port map (
            O => \N__23900\,
            I => \N__23894\
        );

    \I__2696\ : Span4Mux_h
    port map (
            O => \N__23897\,
            I => \N__23891\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__23894\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__23891\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__2693\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23883\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__23883\,
            I => \N__23879\
        );

    \I__2691\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23876\
        );

    \I__2690\ : Span4Mux_v
    port map (
            O => \N__23879\,
            I => \N__23873\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__23876\,
            I => \N__23870\
        );

    \I__2688\ : Span4Mux_v
    port map (
            O => \N__23873\,
            I => \N__23865\
        );

    \I__2687\ : Span4Mux_s3_h
    port map (
            O => \N__23870\,
            I => \N__23865\
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__23865\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__2685\ : InMux
    port map (
            O => \N__23862\,
            I => \N__23859\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__23859\,
            I => \N__23856\
        );

    \I__2683\ : Span4Mux_v
    port map (
            O => \N__23856\,
            I => \N__23852\
        );

    \I__2682\ : InMux
    port map (
            O => \N__23855\,
            I => \N__23849\
        );

    \I__2681\ : Span4Mux_v
    port map (
            O => \N__23852\,
            I => \N__23846\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__23849\,
            I => \N__23843\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__23846\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__2678\ : Odrv12
    port map (
            O => \N__23843\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__2677\ : InMux
    port map (
            O => \N__23838\,
            I => \N__23834\
        );

    \I__2676\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23831\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__23834\,
            I => \N__23828\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__23831\,
            I => \N__23825\
        );

    \I__2673\ : Span4Mux_h
    port map (
            O => \N__23828\,
            I => \N__23822\
        );

    \I__2672\ : Span4Mux_v
    port map (
            O => \N__23825\,
            I => \N__23819\
        );

    \I__2671\ : Span4Mux_v
    port map (
            O => \N__23822\,
            I => \N__23816\
        );

    \I__2670\ : Span4Mux_h
    port map (
            O => \N__23819\,
            I => \N__23813\
        );

    \I__2669\ : Odrv4
    port map (
            O => \N__23816\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__23813\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__2667\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23804\
        );

    \I__2666\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23801\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__23804\,
            I => \N__23798\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__23801\,
            I => \N__23795\
        );

    \I__2663\ : Span4Mux_h
    port map (
            O => \N__23798\,
            I => \N__23792\
        );

    \I__2662\ : Span4Mux_v
    port map (
            O => \N__23795\,
            I => \N__23789\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__23792\,
            I => \N__23786\
        );

    \I__2660\ : Span4Mux_h
    port map (
            O => \N__23789\,
            I => \N__23783\
        );

    \I__2659\ : Odrv4
    port map (
            O => \N__23786\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__23783\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__2657\ : InMux
    port map (
            O => \N__23778\,
            I => \N__23774\
        );

    \I__2656\ : InMux
    port map (
            O => \N__23777\,
            I => \N__23771\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__23774\,
            I => \N__23768\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__23771\,
            I => \N__23765\
        );

    \I__2653\ : Span4Mux_v
    port map (
            O => \N__23768\,
            I => \N__23762\
        );

    \I__2652\ : Span4Mux_v
    port map (
            O => \N__23765\,
            I => \N__23759\
        );

    \I__2651\ : Span4Mux_v
    port map (
            O => \N__23762\,
            I => \N__23756\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__23759\,
            I => \N__23753\
        );

    \I__2649\ : Odrv4
    port map (
            O => \N__23756\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__2648\ : Odrv4
    port map (
            O => \N__23753\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__2647\ : InMux
    port map (
            O => \N__23748\,
            I => \N__23745\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__23745\,
            I => \N__23742\
        );

    \I__2645\ : Span4Mux_v
    port map (
            O => \N__23742\,
            I => \N__23738\
        );

    \I__2644\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23735\
        );

    \I__2643\ : Sp12to4
    port map (
            O => \N__23738\,
            I => \N__23730\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__23735\,
            I => \N__23730\
        );

    \I__2641\ : Span12Mux_s5_h
    port map (
            O => \N__23730\,
            I => \N__23727\
        );

    \I__2640\ : Odrv12
    port map (
            O => \N__23727\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__2639\ : InMux
    port map (
            O => \N__23724\,
            I => \N__23720\
        );

    \I__2638\ : InMux
    port map (
            O => \N__23723\,
            I => \N__23717\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__23720\,
            I => \N__23714\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__23717\,
            I => \N__23711\
        );

    \I__2635\ : Span4Mux_h
    port map (
            O => \N__23714\,
            I => \N__23708\
        );

    \I__2634\ : Span12Mux_s5_h
    port map (
            O => \N__23711\,
            I => \N__23705\
        );

    \I__2633\ : Odrv4
    port map (
            O => \N__23708\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__2632\ : Odrv12
    port map (
            O => \N__23705\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__2631\ : InMux
    port map (
            O => \N__23700\,
            I => \N__23697\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__23697\,
            I => \N__23694\
        );

    \I__2629\ : Span4Mux_h
    port map (
            O => \N__23694\,
            I => \N__23691\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__23691\,
            I => \current_shift_inst.control_input_axb_16\
        );

    \I__2627\ : InMux
    port map (
            O => \N__23688\,
            I => \N__23685\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__23685\,
            I => \N__23682\
        );

    \I__2625\ : Span4Mux_v
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__2624\ : Span4Mux_h
    port map (
            O => \N__23679\,
            I => \N__23676\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__23676\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__2622\ : InMux
    port map (
            O => \N__23673\,
            I => \N__23670\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__23670\,
            I => \N__23666\
        );

    \I__2620\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23663\
        );

    \I__2619\ : Span4Mux_v
    port map (
            O => \N__23666\,
            I => \N__23658\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__23663\,
            I => \N__23658\
        );

    \I__2617\ : Span4Mux_h
    port map (
            O => \N__23658\,
            I => \N__23655\
        );

    \I__2616\ : Span4Mux_v
    port map (
            O => \N__23655\,
            I => \N__23652\
        );

    \I__2615\ : Odrv4
    port map (
            O => \N__23652\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__2614\ : InMux
    port map (
            O => \N__23649\,
            I => \N__23646\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__23646\,
            I => \N__23643\
        );

    \I__2612\ : Span4Mux_h
    port map (
            O => \N__23643\,
            I => \N__23640\
        );

    \I__2611\ : Span4Mux_v
    port map (
            O => \N__23640\,
            I => \N__23637\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__23637\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__2609\ : InMux
    port map (
            O => \N__23634\,
            I => \N__23631\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__23631\,
            I => \N__23628\
        );

    \I__2607\ : Span12Mux_s7_h
    port map (
            O => \N__23628\,
            I => \N__23625\
        );

    \I__2606\ : Odrv12
    port map (
            O => \N__23625\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__2605\ : InMux
    port map (
            O => \N__23622\,
            I => \N__23619\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__23619\,
            I => \N__23615\
        );

    \I__2603\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23612\
        );

    \I__2602\ : Span4Mux_s1_h
    port map (
            O => \N__23615\,
            I => \N__23609\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__23612\,
            I => \N__23606\
        );

    \I__2600\ : Span4Mux_h
    port map (
            O => \N__23609\,
            I => \N__23603\
        );

    \I__2599\ : Odrv4
    port map (
            O => \N__23606\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__23603\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__2597\ : InMux
    port map (
            O => \N__23598\,
            I => \N__23595\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__23595\,
            I => \N__23592\
        );

    \I__2595\ : Span4Mux_h
    port map (
            O => \N__23592\,
            I => \N__23589\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__23589\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__2593\ : InMux
    port map (
            O => \N__23586\,
            I => \N__23583\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__23583\,
            I => \N__23580\
        );

    \I__2591\ : Span4Mux_h
    port map (
            O => \N__23580\,
            I => \N__23577\
        );

    \I__2590\ : Odrv4
    port map (
            O => \N__23577\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__2589\ : InMux
    port map (
            O => \N__23574\,
            I => \N__23571\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__23571\,
            I => \N__23568\
        );

    \I__2587\ : Span4Mux_h
    port map (
            O => \N__23568\,
            I => \N__23565\
        );

    \I__2586\ : Odrv4
    port map (
            O => \N__23565\,
            I => \current_shift_inst.control_input_axb_14\
        );

    \I__2585\ : InMux
    port map (
            O => \N__23562\,
            I => \N__23559\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__23559\,
            I => \N__23556\
        );

    \I__2583\ : Odrv12
    port map (
            O => \N__23556\,
            I => \current_shift_inst.control_input_axb_26\
        );

    \I__2582\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23550\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__23550\,
            I => \N__23547\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__23547\,
            I => \N__23544\
        );

    \I__2579\ : Odrv4
    port map (
            O => \N__23544\,
            I => \current_shift_inst.control_input_axb_21\
        );

    \I__2578\ : InMux
    port map (
            O => \N__23541\,
            I => \N__23538\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__23538\,
            I => \N__23535\
        );

    \I__2576\ : Span4Mux_h
    port map (
            O => \N__23535\,
            I => \N__23532\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__23532\,
            I => \current_shift_inst.control_input_axb_17\
        );

    \I__2574\ : InMux
    port map (
            O => \N__23529\,
            I => \N__23526\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__23526\,
            I => \N__23523\
        );

    \I__2572\ : Span4Mux_h
    port map (
            O => \N__23523\,
            I => \N__23520\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__23520\,
            I => \current_shift_inst.control_input_axb_15\
        );

    \I__2570\ : InMux
    port map (
            O => \N__23517\,
            I => \N__23513\
        );

    \I__2569\ : InMux
    port map (
            O => \N__23516\,
            I => \N__23510\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__23513\,
            I => \N__23507\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__23510\,
            I => \N__23504\
        );

    \I__2566\ : Span4Mux_s1_h
    port map (
            O => \N__23507\,
            I => \N__23501\
        );

    \I__2565\ : Span4Mux_v
    port map (
            O => \N__23504\,
            I => \N__23498\
        );

    \I__2564\ : Span4Mux_h
    port map (
            O => \N__23501\,
            I => \N__23495\
        );

    \I__2563\ : Odrv4
    port map (
            O => \N__23498\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__2562\ : Odrv4
    port map (
            O => \N__23495\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__2561\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23486\
        );

    \I__2560\ : InMux
    port map (
            O => \N__23489\,
            I => \N__23483\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__23486\,
            I => \N__23480\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__23483\,
            I => \N__23477\
        );

    \I__2557\ : Span4Mux_v
    port map (
            O => \N__23480\,
            I => \N__23474\
        );

    \I__2556\ : Span4Mux_v
    port map (
            O => \N__23477\,
            I => \N__23471\
        );

    \I__2555\ : Span4Mux_h
    port map (
            O => \N__23474\,
            I => \N__23468\
        );

    \I__2554\ : Odrv4
    port map (
            O => \N__23471\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__23468\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__2552\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23460\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__23460\,
            I => \N__23456\
        );

    \I__2550\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23453\
        );

    \I__2549\ : Span4Mux_v
    port map (
            O => \N__23456\,
            I => \N__23450\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__23453\,
            I => \N__23447\
        );

    \I__2547\ : Span4Mux_h
    port map (
            O => \N__23450\,
            I => \N__23444\
        );

    \I__2546\ : Odrv12
    port map (
            O => \N__23447\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__2545\ : Odrv4
    port map (
            O => \N__23444\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__2544\ : InMux
    port map (
            O => \N__23439\,
            I => \N__23436\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__23436\,
            I => \N__23432\
        );

    \I__2542\ : InMux
    port map (
            O => \N__23435\,
            I => \N__23429\
        );

    \I__2541\ : Span4Mux_v
    port map (
            O => \N__23432\,
            I => \N__23426\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__23429\,
            I => \N__23423\
        );

    \I__2539\ : Span4Mux_h
    port map (
            O => \N__23426\,
            I => \N__23420\
        );

    \I__2538\ : Odrv12
    port map (
            O => \N__23423\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__23420\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__2536\ : InMux
    port map (
            O => \N__23415\,
            I => \N__23412\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__23412\,
            I => \N__23409\
        );

    \I__2534\ : Odrv12
    port map (
            O => \N__23409\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_31\
        );

    \I__2533\ : InMux
    port map (
            O => \N__23406\,
            I => \N__23403\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__23403\,
            I => \N__23400\
        );

    \I__2531\ : Span4Mux_s1_h
    port map (
            O => \N__23400\,
            I => \N__23396\
        );

    \I__2530\ : InMux
    port map (
            O => \N__23399\,
            I => \N__23393\
        );

    \I__2529\ : Span4Mux_v
    port map (
            O => \N__23396\,
            I => \N__23390\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__23393\,
            I => \N__23387\
        );

    \I__2527\ : Span4Mux_h
    port map (
            O => \N__23390\,
            I => \N__23384\
        );

    \I__2526\ : Odrv12
    port map (
            O => \N__23387\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__23384\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__2524\ : InMux
    port map (
            O => \N__23379\,
            I => \N__23375\
        );

    \I__2523\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23372\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__23375\,
            I => \N__23369\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__23372\,
            I => \N__23366\
        );

    \I__2520\ : Span12Mux_v
    port map (
            O => \N__23369\,
            I => \N__23363\
        );

    \I__2519\ : Odrv12
    port map (
            O => \N__23366\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__2518\ : Odrv12
    port map (
            O => \N__23363\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__2517\ : InMux
    port map (
            O => \N__23358\,
            I => \N__23355\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__23355\,
            I => \N__23351\
        );

    \I__2515\ : InMux
    port map (
            O => \N__23354\,
            I => \N__23348\
        );

    \I__2514\ : Span4Mux_v
    port map (
            O => \N__23351\,
            I => \N__23345\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__23348\,
            I => \N__23342\
        );

    \I__2512\ : Span4Mux_v
    port map (
            O => \N__23345\,
            I => \N__23339\
        );

    \I__2511\ : Span12Mux_s10_v
    port map (
            O => \N__23342\,
            I => \N__23336\
        );

    \I__2510\ : Span4Mux_h
    port map (
            O => \N__23339\,
            I => \N__23333\
        );

    \I__2509\ : Odrv12
    port map (
            O => \N__23336\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__23333\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__2507\ : ClkMux
    port map (
            O => \N__23328\,
            I => \N__23325\
        );

    \I__2506\ : GlobalMux
    port map (
            O => \N__23325\,
            I => \N__23322\
        );

    \I__2505\ : gio2CtrlBuf
    port map (
            O => \N__23322\,
            I => delay_hc_input_c_g
        );

    \I__2504\ : InMux
    port map (
            O => \N__23319\,
            I => \N__23315\
        );

    \I__2503\ : InMux
    port map (
            O => \N__23318\,
            I => \N__23312\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23309\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__23312\,
            I => \N__23306\
        );

    \I__2500\ : Span4Mux_s2_h
    port map (
            O => \N__23309\,
            I => \N__23303\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__23306\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__23303\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__2497\ : InMux
    port map (
            O => \N__23298\,
            I => \N__23294\
        );

    \I__2496\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23291\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__23294\,
            I => \N__23288\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__23291\,
            I => \N__23285\
        );

    \I__2493\ : Odrv12
    port map (
            O => \N__23288\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__2492\ : Odrv12
    port map (
            O => \N__23285\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__2491\ : InMux
    port map (
            O => \N__23280\,
            I => \N__23276\
        );

    \I__2490\ : InMux
    port map (
            O => \N__23279\,
            I => \N__23273\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__23276\,
            I => \N__23270\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__23273\,
            I => \N__23267\
        );

    \I__2487\ : Span4Mux_s3_h
    port map (
            O => \N__23270\,
            I => \N__23264\
        );

    \I__2486\ : Odrv12
    port map (
            O => \N__23267\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__2485\ : Odrv4
    port map (
            O => \N__23264\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__2484\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23256\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__23256\,
            I => \N__23252\
        );

    \I__2482\ : InMux
    port map (
            O => \N__23255\,
            I => \N__23249\
        );

    \I__2481\ : Span4Mux_v
    port map (
            O => \N__23252\,
            I => \N__23246\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__23249\,
            I => \N__23243\
        );

    \I__2479\ : Span4Mux_h
    port map (
            O => \N__23246\,
            I => \N__23240\
        );

    \I__2478\ : Odrv4
    port map (
            O => \N__23243\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__23240\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__2476\ : InMux
    port map (
            O => \N__23235\,
            I => \N__23232\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__23232\,
            I => \N__23228\
        );

    \I__2474\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23225\
        );

    \I__2473\ : Span4Mux_v
    port map (
            O => \N__23228\,
            I => \N__23222\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__23225\,
            I => \N__23219\
        );

    \I__2471\ : Span4Mux_h
    port map (
            O => \N__23222\,
            I => \N__23216\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__23219\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__2469\ : Odrv4
    port map (
            O => \N__23216\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__2468\ : InMux
    port map (
            O => \N__23211\,
            I => \N__23208\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__23208\,
            I => \N__23204\
        );

    \I__2466\ : InMux
    port map (
            O => \N__23207\,
            I => \N__23201\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__23204\,
            I => \N__23198\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__23201\,
            I => \N__23195\
        );

    \I__2463\ : Span4Mux_h
    port map (
            O => \N__23198\,
            I => \N__23192\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__23195\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_27\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__23192\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_27\
        );

    \I__2460\ : InMux
    port map (
            O => \N__23187\,
            I => \N__23184\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__23184\,
            I => \N__23180\
        );

    \I__2458\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23177\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__23180\,
            I => \N__23174\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__23177\,
            I => \N__23171\
        );

    \I__2455\ : Span4Mux_h
    port map (
            O => \N__23174\,
            I => \N__23168\
        );

    \I__2454\ : Odrv12
    port map (
            O => \N__23171\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__23168\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__2452\ : InMux
    port map (
            O => \N__23163\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_24\
        );

    \I__2451\ : InMux
    port map (
            O => \N__23160\,
            I => \N__23157\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__23157\,
            I => \N__23154\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__23154\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\
        );

    \I__2448\ : InMux
    port map (
            O => \N__23151\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_25\
        );

    \I__2447\ : InMux
    port map (
            O => \N__23148\,
            I => \N__23145\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__23145\,
            I => \N__23142\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__23142\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\
        );

    \I__2444\ : InMux
    port map (
            O => \N__23139\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_26\
        );

    \I__2443\ : InMux
    port map (
            O => \N__23136\,
            I => \N__23133\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__23133\,
            I => \N__23130\
        );

    \I__2441\ : Odrv12
    port map (
            O => \N__23130\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\
        );

    \I__2440\ : InMux
    port map (
            O => \N__23127\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_27\
        );

    \I__2439\ : InMux
    port map (
            O => \N__23124\,
            I => \N__23121\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__23121\,
            I => \N__23118\
        );

    \I__2437\ : Odrv12
    port map (
            O => \N__23118\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\
        );

    \I__2436\ : InMux
    port map (
            O => \N__23115\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_28\
        );

    \I__2435\ : InMux
    port map (
            O => \N__23112\,
            I => \N__23109\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__23109\,
            I => \N__23106\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__23106\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\
        );

    \I__2432\ : InMux
    port map (
            O => \N__23103\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_29\
        );

    \I__2431\ : InMux
    port map (
            O => \N__23100\,
            I => \N__23097\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__23097\,
            I => \N__23094\
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__23094\,
            I => \current_shift_inst.control_input_31\
        );

    \I__2428\ : InMux
    port map (
            O => \N__23091\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_30\
        );

    \I__2427\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23084\
        );

    \I__2426\ : InMux
    port map (
            O => \N__23087\,
            I => \N__23081\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__23084\,
            I => \N__23078\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__23081\,
            I => \N__23075\
        );

    \I__2423\ : Span4Mux_s1_h
    port map (
            O => \N__23078\,
            I => \N__23072\
        );

    \I__2422\ : Span4Mux_v
    port map (
            O => \N__23075\,
            I => \N__23067\
        );

    \I__2421\ : Span4Mux_h
    port map (
            O => \N__23072\,
            I => \N__23067\
        );

    \I__2420\ : Odrv4
    port map (
            O => \N__23067\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__2419\ : InMux
    port map (
            O => \N__23064\,
            I => \N__23061\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__23061\,
            I => \N__23057\
        );

    \I__2417\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23054\
        );

    \I__2416\ : Span4Mux_v
    port map (
            O => \N__23057\,
            I => \N__23051\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__23054\,
            I => \N__23048\
        );

    \I__2414\ : Span4Mux_h
    port map (
            O => \N__23051\,
            I => \N__23045\
        );

    \I__2413\ : Odrv4
    port map (
            O => \N__23048\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__2412\ : Odrv4
    port map (
            O => \N__23045\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__2411\ : InMux
    port map (
            O => \N__23040\,
            I => \N__23037\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__23037\,
            I => \N__23034\
        );

    \I__2409\ : Odrv4
    port map (
            O => \N__23034\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\
        );

    \I__2408\ : InMux
    port map (
            O => \N__23031\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_16\
        );

    \I__2407\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23025\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__23025\,
            I => \N__23022\
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__23022\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\
        );

    \I__2404\ : InMux
    port map (
            O => \N__23019\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_17\
        );

    \I__2403\ : InMux
    port map (
            O => \N__23016\,
            I => \N__23013\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__23013\,
            I => \N__23010\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__23010\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\
        );

    \I__2400\ : InMux
    port map (
            O => \N__23007\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_18\
        );

    \I__2399\ : InMux
    port map (
            O => \N__23004\,
            I => \N__23001\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__23001\,
            I => \N__22998\
        );

    \I__2397\ : Odrv12
    port map (
            O => \N__22998\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\
        );

    \I__2396\ : InMux
    port map (
            O => \N__22995\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_19\
        );

    \I__2395\ : InMux
    port map (
            O => \N__22992\,
            I => \N__22989\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__22989\,
            I => \N__22986\
        );

    \I__2393\ : Odrv12
    port map (
            O => \N__22986\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\
        );

    \I__2392\ : InMux
    port map (
            O => \N__22983\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_20\
        );

    \I__2391\ : InMux
    port map (
            O => \N__22980\,
            I => \N__22977\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__22977\,
            I => \N__22974\
        );

    \I__2389\ : Odrv12
    port map (
            O => \N__22974\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\
        );

    \I__2388\ : InMux
    port map (
            O => \N__22971\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_21\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__22968\,
            I => \N__22965\
        );

    \I__2386\ : InMux
    port map (
            O => \N__22965\,
            I => \N__22962\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__22962\,
            I => \N__22959\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__22959\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\
        );

    \I__2383\ : InMux
    port map (
            O => \N__22956\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_22\
        );

    \I__2382\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22950\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__22950\,
            I => \N__22947\
        );

    \I__2380\ : Odrv4
    port map (
            O => \N__22947\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\
        );

    \I__2379\ : InMux
    port map (
            O => \N__22944\,
            I => \bfn_5_14_0_\
        );

    \I__2378\ : InMux
    port map (
            O => \N__22941\,
            I => \N__22938\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__22938\,
            I => \N__22935\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__22935\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\
        );

    \I__2375\ : InMux
    port map (
            O => \N__22932\,
            I => \N__22929\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__22929\,
            I => \N__22926\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__22926\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__2372\ : InMux
    port map (
            O => \N__22923\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__2371\ : InMux
    port map (
            O => \N__22920\,
            I => \N__22917\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__22917\,
            I => \N__22914\
        );

    \I__2369\ : Odrv4
    port map (
            O => \N__22914\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__2368\ : InMux
    port map (
            O => \N__22911\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__2367\ : CascadeMux
    port map (
            O => \N__22908\,
            I => \N__22905\
        );

    \I__2366\ : InMux
    port map (
            O => \N__22905\,
            I => \N__22902\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__22902\,
            I => \N__22899\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__22899\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__2363\ : InMux
    port map (
            O => \N__22896\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__2362\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22890\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__22890\,
            I => \N__22887\
        );

    \I__2360\ : Odrv12
    port map (
            O => \N__22887\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__2359\ : InMux
    port map (
            O => \N__22884\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__2358\ : InMux
    port map (
            O => \N__22881\,
            I => \N__22878\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__22878\,
            I => \N__22875\
        );

    \I__2356\ : Odrv12
    port map (
            O => \N__22875\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__2355\ : InMux
    port map (
            O => \N__22872\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__2354\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22866\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__22866\,
            I => \N__22863\
        );

    \I__2352\ : Odrv12
    port map (
            O => \N__22863\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\
        );

    \I__2351\ : InMux
    port map (
            O => \N__22860\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__2350\ : InMux
    port map (
            O => \N__22857\,
            I => \N__22854\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__22854\,
            I => \N__22851\
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__22851\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\
        );

    \I__2347\ : InMux
    port map (
            O => \N__22848\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_14\
        );

    \I__2346\ : InMux
    port map (
            O => \N__22845\,
            I => \N__22842\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__22842\,
            I => \N__22839\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__22839\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\
        );

    \I__2343\ : InMux
    port map (
            O => \N__22836\,
            I => \bfn_5_13_0_\
        );

    \I__2342\ : InMux
    port map (
            O => \N__22833\,
            I => \N__22830\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__22830\,
            I => \N__22827\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__22827\,
            I => \current_shift_inst.control_input_1\
        );

    \I__2339\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22821\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__22821\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__2337\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22815\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__22815\,
            I => \N__22812\
        );

    \I__2335\ : Odrv4
    port map (
            O => \N__22812\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__2334\ : InMux
    port map (
            O => \N__22809\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__22806\,
            I => \N__22803\
        );

    \I__2332\ : InMux
    port map (
            O => \N__22803\,
            I => \N__22800\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__22800\,
            I => \N__22797\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__22797\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__2329\ : InMux
    port map (
            O => \N__22794\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__2328\ : InMux
    port map (
            O => \N__22791\,
            I => \N__22788\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__22788\,
            I => \N__22785\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__22785\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__2325\ : InMux
    port map (
            O => \N__22782\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__2324\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22776\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__22776\,
            I => \N__22773\
        );

    \I__2322\ : Odrv12
    port map (
            O => \N__22773\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__2321\ : InMux
    port map (
            O => \N__22770\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__2320\ : InMux
    port map (
            O => \N__22767\,
            I => \N__22764\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__22764\,
            I => \N__22761\
        );

    \I__2318\ : Odrv12
    port map (
            O => \N__22761\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__2317\ : InMux
    port map (
            O => \N__22758\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__2316\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22752\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__22752\,
            I => \N__22749\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__22749\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__2313\ : InMux
    port map (
            O => \N__22746\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__2312\ : InMux
    port map (
            O => \N__22743\,
            I => \N__22740\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__22740\,
            I => \N__22737\
        );

    \I__2310\ : Odrv12
    port map (
            O => \N__22737\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__2309\ : InMux
    port map (
            O => \N__22734\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__2308\ : InMux
    port map (
            O => \N__22731\,
            I => \N__22728\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__22728\,
            I => \N__22725\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__22725\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__2305\ : InMux
    port map (
            O => \N__22722\,
            I => \bfn_5_12_0_\
        );

    \I__2304\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22716\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__22716\,
            I => \current_shift_inst.control_input_axb_23\
        );

    \I__2302\ : InMux
    port map (
            O => \N__22713\,
            I => \N__22710\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__22710\,
            I => \current_shift_inst.control_input_axb_25\
        );

    \I__2300\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22704\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__22704\,
            I => \N__22701\
        );

    \I__2298\ : Span4Mux_h
    port map (
            O => \N__22701\,
            I => \N__22698\
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__22698\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__2296\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22692\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__22692\,
            I => \current_shift_inst.control_input_axb_29\
        );

    \I__2294\ : CascadeMux
    port map (
            O => \N__22689\,
            I => \current_shift_inst.PI_CTRL.N_46_16_cascade_\
        );

    \I__2293\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22683\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__22683\,
            I => \N__22680\
        );

    \I__2291\ : Odrv12
    port map (
            O => \N__22680\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\
        );

    \I__2290\ : InMux
    port map (
            O => \N__22677\,
            I => \N__22674\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__22674\,
            I => \N__22670\
        );

    \I__2288\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22667\
        );

    \I__2287\ : Span4Mux_v
    port map (
            O => \N__22670\,
            I => \N__22664\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__22667\,
            I => \N__22661\
        );

    \I__2285\ : Span4Mux_v
    port map (
            O => \N__22664\,
            I => \N__22656\
        );

    \I__2284\ : Span4Mux_h
    port map (
            O => \N__22661\,
            I => \N__22656\
        );

    \I__2283\ : Odrv4
    port map (
            O => \N__22656\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__22653\,
            I => \N__22643\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__22652\,
            I => \N__22640\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__22651\,
            I => \N__22637\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__22650\,
            I => \N__22634\
        );

    \I__2278\ : CEMux
    port map (
            O => \N__22649\,
            I => \N__22629\
        );

    \I__2277\ : InMux
    port map (
            O => \N__22648\,
            I => \N__22617\
        );

    \I__2276\ : InMux
    port map (
            O => \N__22647\,
            I => \N__22614\
        );

    \I__2275\ : InMux
    port map (
            O => \N__22646\,
            I => \N__22611\
        );

    \I__2274\ : InMux
    port map (
            O => \N__22643\,
            I => \N__22598\
        );

    \I__2273\ : InMux
    port map (
            O => \N__22640\,
            I => \N__22598\
        );

    \I__2272\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22598\
        );

    \I__2271\ : InMux
    port map (
            O => \N__22634\,
            I => \N__22598\
        );

    \I__2270\ : InMux
    port map (
            O => \N__22633\,
            I => \N__22598\
        );

    \I__2269\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22598\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__22629\,
            I => \N__22592\
        );

    \I__2267\ : InMux
    port map (
            O => \N__22628\,
            I => \N__22587\
        );

    \I__2266\ : InMux
    port map (
            O => \N__22627\,
            I => \N__22587\
        );

    \I__2265\ : InMux
    port map (
            O => \N__22626\,
            I => \N__22580\
        );

    \I__2264\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22580\
        );

    \I__2263\ : InMux
    port map (
            O => \N__22624\,
            I => \N__22580\
        );

    \I__2262\ : InMux
    port map (
            O => \N__22623\,
            I => \N__22573\
        );

    \I__2261\ : InMux
    port map (
            O => \N__22622\,
            I => \N__22573\
        );

    \I__2260\ : InMux
    port map (
            O => \N__22621\,
            I => \N__22573\
        );

    \I__2259\ : InMux
    port map (
            O => \N__22620\,
            I => \N__22570\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__22617\,
            I => \N__22567\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__22614\,
            I => \N__22564\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__22611\,
            I => \N__22559\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__22598\,
            I => \N__22559\
        );

    \I__2254\ : InMux
    port map (
            O => \N__22597\,
            I => \N__22545\
        );

    \I__2253\ : InMux
    port map (
            O => \N__22596\,
            I => \N__22545\
        );

    \I__2252\ : InMux
    port map (
            O => \N__22595\,
            I => \N__22542\
        );

    \I__2251\ : Span4Mux_h
    port map (
            O => \N__22592\,
            I => \N__22533\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__22587\,
            I => \N__22533\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__22580\,
            I => \N__22533\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__22573\,
            I => \N__22533\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__22570\,
            I => \N__22528\
        );

    \I__2246\ : Span4Mux_h
    port map (
            O => \N__22567\,
            I => \N__22528\
        );

    \I__2245\ : Span4Mux_h
    port map (
            O => \N__22564\,
            I => \N__22523\
        );

    \I__2244\ : Span4Mux_h
    port map (
            O => \N__22559\,
            I => \N__22523\
        );

    \I__2243\ : InMux
    port map (
            O => \N__22558\,
            I => \N__22520\
        );

    \I__2242\ : InMux
    port map (
            O => \N__22557\,
            I => \N__22511\
        );

    \I__2241\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22511\
        );

    \I__2240\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22511\
        );

    \I__2239\ : InMux
    port map (
            O => \N__22554\,
            I => \N__22511\
        );

    \I__2238\ : InMux
    port map (
            O => \N__22553\,
            I => \N__22502\
        );

    \I__2237\ : InMux
    port map (
            O => \N__22552\,
            I => \N__22502\
        );

    \I__2236\ : InMux
    port map (
            O => \N__22551\,
            I => \N__22502\
        );

    \I__2235\ : InMux
    port map (
            O => \N__22550\,
            I => \N__22502\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__22545\,
            I => \N__22499\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__22542\,
            I => \N__22494\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__22533\,
            I => \N__22494\
        );

    \I__2231\ : Span4Mux_v
    port map (
            O => \N__22528\,
            I => \N__22491\
        );

    \I__2230\ : Span4Mux_v
    port map (
            O => \N__22523\,
            I => \N__22488\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__22520\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__22511\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__22502\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__2226\ : Odrv12
    port map (
            O => \N__22499\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__2225\ : Odrv4
    port map (
            O => \N__22494\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__22491\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__22488\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__2222\ : InMux
    port map (
            O => \N__22473\,
            I => \N__22470\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__22470\,
            I => \N__22467\
        );

    \I__2220\ : Span4Mux_v
    port map (
            O => \N__22467\,
            I => \N__22464\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__22464\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__2218\ : InMux
    port map (
            O => \N__22461\,
            I => \N__22458\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__22458\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__2216\ : InMux
    port map (
            O => \N__22455\,
            I => \N__22452\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__22452\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__2214\ : InMux
    port map (
            O => \N__22449\,
            I => \N__22446\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__22446\,
            I => \current_shift_inst.control_input_axb_13\
        );

    \I__2212\ : InMux
    port map (
            O => \N__22443\,
            I => \N__22440\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__22440\,
            I => \current_shift_inst.control_input_axb_18\
        );

    \I__2210\ : InMux
    port map (
            O => \N__22437\,
            I => \N__22434\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__22434\,
            I => \current_shift_inst.control_input_axb_20\
        );

    \I__2208\ : InMux
    port map (
            O => \N__22431\,
            I => \N__22428\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__22428\,
            I => \N__22425\
        );

    \I__2206\ : Odrv12
    port map (
            O => \N__22425\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\
        );

    \I__2205\ : InMux
    port map (
            O => \N__22422\,
            I => \N__22419\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__22419\,
            I => \N__22416\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__22416\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__2202\ : InMux
    port map (
            O => \N__22413\,
            I => \N__22410\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__22410\,
            I => \current_shift_inst.control_input_axb_27\
        );

    \I__2200\ : InMux
    port map (
            O => \N__22407\,
            I => \N__22404\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__22404\,
            I => \current_shift_inst.control_input_axb_22\
        );

    \I__2198\ : InMux
    port map (
            O => \N__22401\,
            I => \N__22398\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__22398\,
            I => \current_shift_inst.control_input_axb_24\
        );

    \I__2196\ : InMux
    port map (
            O => \N__22395\,
            I => \N__22392\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__22392\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__2194\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22386\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__22386\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\
        );

    \I__2192\ : InMux
    port map (
            O => \N__22383\,
            I => \N__22380\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__22380\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\
        );

    \I__2190\ : InMux
    port map (
            O => \N__22377\,
            I => \N__22374\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__22374\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__2188\ : InMux
    port map (
            O => \N__22371\,
            I => \N__22368\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__22368\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__2186\ : InMux
    port map (
            O => \N__22365\,
            I => \N__22362\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__22362\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__2184\ : InMux
    port map (
            O => \N__22359\,
            I => \N__22356\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__22356\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__2182\ : InMux
    port map (
            O => \N__22353\,
            I => \N__22350\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__22350\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__22347\,
            I => \N__22344\
        );

    \I__2179\ : InMux
    port map (
            O => \N__22344\,
            I => \N__22341\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__22341\,
            I => \N__22338\
        );

    \I__2177\ : Odrv4
    port map (
            O => \N__22338\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__22335\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_\
        );

    \I__2175\ : InMux
    port map (
            O => \N__22332\,
            I => \N__22329\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__22329\,
            I => \current_shift_inst.PI_CTRL.N_77\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__22326\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\
        );

    \I__2172\ : CascadeMux
    port map (
            O => \N__22323\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\
        );

    \I__2171\ : InMux
    port map (
            O => \N__22320\,
            I => \N__22317\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__22317\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__2169\ : InMux
    port map (
            O => \N__22314\,
            I => \N__22311\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__22311\,
            I => \N__22308\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__22308\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2166\ : InMux
    port map (
            O => \N__22305\,
            I => \N__22302\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__22302\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\
        );

    \I__2164\ : InMux
    port map (
            O => \N__22299\,
            I => \N__22296\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__22296\,
            I => \N__22293\
        );

    \I__2162\ : Odrv4
    port map (
            O => \N__22293\,
            I => \current_shift_inst.PI_CTRL.N_46_21\
        );

    \I__2161\ : InMux
    port map (
            O => \N__22290\,
            I => \N__22287\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__22287\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__2159\ : InMux
    port map (
            O => \N__22284\,
            I => \current_shift_inst.control_input_cry_26\
        );

    \I__2158\ : InMux
    port map (
            O => \N__22281\,
            I => \current_shift_inst.control_input_cry_27\
        );

    \I__2157\ : InMux
    port map (
            O => \N__22278\,
            I => \current_shift_inst.control_input_cry_28\
        );

    \I__2156\ : InMux
    port map (
            O => \N__22275\,
            I => \current_shift_inst.control_input_cry_29\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__22272\,
            I => \current_shift_inst.control_input_31_cascade_\
        );

    \I__2154\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22266\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__22266\,
            I => \N__22263\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__22263\,
            I => \N__22260\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__22260\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__2150\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22254\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__22254\,
            I => \N__22251\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__22251\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__22248\,
            I => \current_shift_inst.PI_CTRL.N_44_cascade_\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__22245\,
            I => \N__22240\
        );

    \I__2145\ : InMux
    port map (
            O => \N__22244\,
            I => \N__22237\
        );

    \I__2144\ : InMux
    port map (
            O => \N__22243\,
            I => \N__22234\
        );

    \I__2143\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22231\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__22237\,
            I => \current_shift_inst.N_1571_i\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__22234\,
            I => \current_shift_inst.N_1571_i\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__22231\,
            I => \current_shift_inst.N_1571_i\
        );

    \I__2139\ : InMux
    port map (
            O => \N__22224\,
            I => \current_shift_inst.control_input_cry_17\
        );

    \I__2138\ : InMux
    port map (
            O => \N__22221\,
            I => \current_shift_inst.control_input_cry_18\
        );

    \I__2137\ : InMux
    port map (
            O => \N__22218\,
            I => \current_shift_inst.control_input_cry_19\
        );

    \I__2136\ : InMux
    port map (
            O => \N__22215\,
            I => \current_shift_inst.control_input_cry_20\
        );

    \I__2135\ : InMux
    port map (
            O => \N__22212\,
            I => \current_shift_inst.control_input_cry_21\
        );

    \I__2134\ : InMux
    port map (
            O => \N__22209\,
            I => \current_shift_inst.control_input_cry_22\
        );

    \I__2133\ : InMux
    port map (
            O => \N__22206\,
            I => \bfn_3_14_0_\
        );

    \I__2132\ : InMux
    port map (
            O => \N__22203\,
            I => \current_shift_inst.control_input_cry_24\
        );

    \I__2131\ : InMux
    port map (
            O => \N__22200\,
            I => \current_shift_inst.control_input_cry_25\
        );

    \I__2130\ : InMux
    port map (
            O => \N__22197\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__2129\ : InMux
    port map (
            O => \N__22194\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__2128\ : InMux
    port map (
            O => \N__22191\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__2127\ : InMux
    port map (
            O => \N__22188\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__2126\ : InMux
    port map (
            O => \N__22185\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__2125\ : InMux
    port map (
            O => \N__22182\,
            I => \current_shift_inst.control_input_cry_13\
        );

    \I__2124\ : InMux
    port map (
            O => \N__22179\,
            I => \current_shift_inst.control_input_cry_14\
        );

    \I__2123\ : InMux
    port map (
            O => \N__22176\,
            I => \bfn_3_13_0_\
        );

    \I__2122\ : InMux
    port map (
            O => \N__22173\,
            I => \current_shift_inst.control_input_cry_16\
        );

    \I__2121\ : InMux
    port map (
            O => \N__22170\,
            I => \N__22167\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__22167\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__2119\ : InMux
    port map (
            O => \N__22164\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__2118\ : InMux
    port map (
            O => \N__22161\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__2117\ : InMux
    port map (
            O => \N__22158\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__2116\ : InMux
    port map (
            O => \N__22155\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__2115\ : InMux
    port map (
            O => \N__22152\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__2114\ : InMux
    port map (
            O => \N__22149\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__2113\ : InMux
    port map (
            O => \N__22146\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__2112\ : InMux
    port map (
            O => \N__22143\,
            I => \bfn_3_12_0_\
        );

    \I__2111\ : InMux
    port map (
            O => \N__22140\,
            I => \N__22137\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__22137\,
            I => \N__22134\
        );

    \I__2109\ : Odrv12
    port map (
            O => \N__22134\,
            I => un8_start_stop
        );

    \I__2108\ : InMux
    port map (
            O => \N__22131\,
            I => \N__22128\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__22128\,
            I => \N__22125\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__22125\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__22122\,
            I => \N__22119\
        );

    \I__2104\ : InMux
    port map (
            O => \N__22119\,
            I => \N__22116\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__22116\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__2102\ : InMux
    port map (
            O => \N__22113\,
            I => \N__22110\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__22110\,
            I => \N__22107\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__22107\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__2099\ : InMux
    port map (
            O => \N__22104\,
            I => \N__22101\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__22101\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__2097\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22095\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__22095\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__2095\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22089\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__22089\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__2093\ : InMux
    port map (
            O => \N__22086\,
            I => \N__22083\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__22083\,
            I => \N__22080\
        );

    \I__2091\ : Odrv4
    port map (
            O => \N__22080\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__2090\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22074\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__22074\,
            I => \N__22071\
        );

    \I__2088\ : Odrv4
    port map (
            O => \N__22071\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__22068\,
            I => \N__22065\
        );

    \I__2086\ : InMux
    port map (
            O => \N__22065\,
            I => \N__22062\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__22062\,
            I => \N__22059\
        );

    \I__2084\ : Span4Mux_v
    port map (
            O => \N__22059\,
            I => \N__22056\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__22056\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\
        );

    \I__2082\ : InMux
    port map (
            O => \N__22053\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__2081\ : InMux
    port map (
            O => \N__22050\,
            I => \N__22047\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__22047\,
            I => \N__22044\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__22044\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__2078\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22038\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__22038\,
            I => \N__22035\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__22035\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__2075\ : InMux
    port map (
            O => \N__22032\,
            I => \N__22029\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__22029\,
            I => \N__22026\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__22026\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__2072\ : InMux
    port map (
            O => \N__22023\,
            I => \N__22020\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__22020\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__2070\ : InMux
    port map (
            O => \N__22017\,
            I => \N__22014\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__22014\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__2068\ : InMux
    port map (
            O => \N__22011\,
            I => \N__22008\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__22008\,
            I => \N__22005\
        );

    \I__2066\ : Odrv4
    port map (
            O => \N__22005\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__2065\ : InMux
    port map (
            O => \N__22002\,
            I => \N__21999\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__21999\,
            I => \N__21996\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__21996\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__2062\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21990\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__21990\,
            I => \N__21987\
        );

    \I__2060\ : Glb2LocalMux
    port map (
            O => \N__21987\,
            I => \N__21984\
        );

    \I__2059\ : GlobalMux
    port map (
            O => \N__21984\,
            I => clk_12mhz
        );

    \I__2058\ : IoInMux
    port map (
            O => \N__21981\,
            I => \N__21978\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__21978\,
            I => \N__21975\
        );

    \I__2056\ : Span4Mux_s0_v
    port map (
            O => \N__21975\,
            I => \N__21972\
        );

    \I__2055\ : Span4Mux_h
    port map (
            O => \N__21972\,
            I => \N__21969\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__21969\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__21966\,
            I => \N__21963\
        );

    \I__2052\ : InMux
    port map (
            O => \N__21963\,
            I => \N__21960\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__21960\,
            I => \N__21957\
        );

    \I__2050\ : Odrv4
    port map (
            O => \N__21957\,
            I => \current_shift_inst.PI_CTRL.integrator_1_23\
        );

    \I__2049\ : InMux
    port map (
            O => \N__21954\,
            I => \N__21951\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__21951\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__2047\ : InMux
    port map (
            O => \N__21948\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__21945\,
            I => \N__21942\
        );

    \I__2045\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21939\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__21939\,
            I => \N__21936\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__21936\,
            I => \current_shift_inst.PI_CTRL.integrator_1_24\
        );

    \I__2042\ : InMux
    port map (
            O => \N__21933\,
            I => \N__21930\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__21930\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__2040\ : InMux
    port map (
            O => \N__21927\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__21924\,
            I => \N__21921\
        );

    \I__2038\ : InMux
    port map (
            O => \N__21921\,
            I => \N__21918\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__21918\,
            I => \N__21915\
        );

    \I__2036\ : Span4Mux_v
    port map (
            O => \N__21915\,
            I => \N__21912\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__21912\,
            I => \current_shift_inst.PI_CTRL.integrator_1_25\
        );

    \I__2034\ : InMux
    port map (
            O => \N__21909\,
            I => \bfn_2_13_0_\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__21906\,
            I => \N__21903\
        );

    \I__2032\ : InMux
    port map (
            O => \N__21903\,
            I => \N__21900\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__21900\,
            I => \N__21897\
        );

    \I__2030\ : Span4Mux_v
    port map (
            O => \N__21897\,
            I => \N__21894\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__21894\,
            I => \current_shift_inst.PI_CTRL.integrator_1_26\
        );

    \I__2028\ : InMux
    port map (
            O => \N__21891\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__21888\,
            I => \N__21885\
        );

    \I__2026\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21882\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__21882\,
            I => \N__21879\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__21879\,
            I => \N__21876\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__21876\,
            I => \current_shift_inst.PI_CTRL.integrator_1_27\
        );

    \I__2022\ : InMux
    port map (
            O => \N__21873\,
            I => \N__21870\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__21870\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__2020\ : InMux
    port map (
            O => \N__21867\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__2019\ : InMux
    port map (
            O => \N__21864\,
            I => \N__21861\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__21861\,
            I => \N__21858\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__21858\,
            I => \current_shift_inst.PI_CTRL.integrator_1_28\
        );

    \I__2016\ : InMux
    port map (
            O => \N__21855\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__21852\,
            I => \N__21849\
        );

    \I__2014\ : InMux
    port map (
            O => \N__21849\,
            I => \N__21846\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__21846\,
            I => \N__21843\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__21843\,
            I => \current_shift_inst.PI_CTRL.integrator_1_29\
        );

    \I__2011\ : InMux
    port map (
            O => \N__21840\,
            I => \N__21837\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__21837\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__2009\ : InMux
    port map (
            O => \N__21834\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__21831\,
            I => \N__21828\
        );

    \I__2007\ : InMux
    port map (
            O => \N__21828\,
            I => \N__21825\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__21825\,
            I => \N__21822\
        );

    \I__2005\ : Span4Mux_v
    port map (
            O => \N__21822\,
            I => \N__21819\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__21819\,
            I => \current_shift_inst.PI_CTRL.integrator_1_30\
        );

    \I__2003\ : InMux
    port map (
            O => \N__21816\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__21813\,
            I => \N__21810\
        );

    \I__2001\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21807\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__21807\,
            I => \N__21804\
        );

    \I__1999\ : Span4Mux_v
    port map (
            O => \N__21804\,
            I => \N__21801\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__21801\,
            I => \current_shift_inst.PI_CTRL.integrator_1_15\
        );

    \I__1997\ : InMux
    port map (
            O => \N__21798\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__21795\,
            I => \N__21792\
        );

    \I__1995\ : InMux
    port map (
            O => \N__21792\,
            I => \N__21789\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__21789\,
            I => \current_shift_inst.PI_CTRL.integrator_1_16\
        );

    \I__1993\ : InMux
    port map (
            O => \N__21786\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__21783\,
            I => \N__21780\
        );

    \I__1991\ : InMux
    port map (
            O => \N__21780\,
            I => \N__21777\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__21777\,
            I => \N__21774\
        );

    \I__1989\ : Span4Mux_v
    port map (
            O => \N__21774\,
            I => \N__21771\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__21771\,
            I => \current_shift_inst.PI_CTRL.integrator_1_17\
        );

    \I__1987\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21765\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__21765\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__1985\ : InMux
    port map (
            O => \N__21762\,
            I => \bfn_2_12_0_\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__21759\,
            I => \N__21756\
        );

    \I__1983\ : InMux
    port map (
            O => \N__21756\,
            I => \N__21753\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__21753\,
            I => \N__21750\
        );

    \I__1981\ : Odrv4
    port map (
            O => \N__21750\,
            I => \current_shift_inst.PI_CTRL.integrator_1_18\
        );

    \I__1980\ : InMux
    port map (
            O => \N__21747\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__21744\,
            I => \N__21741\
        );

    \I__1978\ : InMux
    port map (
            O => \N__21741\,
            I => \N__21738\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__21738\,
            I => \N__21735\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__21735\,
            I => \N__21732\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__21732\,
            I => \current_shift_inst.PI_CTRL.integrator_1_19\
        );

    \I__1974\ : InMux
    port map (
            O => \N__21729\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__1973\ : InMux
    port map (
            O => \N__21726\,
            I => \N__21723\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__21723\,
            I => \N__21720\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__21720\,
            I => \current_shift_inst.PI_CTRL.integrator_1_20\
        );

    \I__1970\ : InMux
    port map (
            O => \N__21717\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__21714\,
            I => \N__21711\
        );

    \I__1968\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21708\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__21708\,
            I => \N__21705\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__21705\,
            I => \current_shift_inst.PI_CTRL.integrator_1_21\
        );

    \I__1965\ : InMux
    port map (
            O => \N__21702\,
            I => \N__21699\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__21699\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__1963\ : InMux
    port map (
            O => \N__21696\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__21693\,
            I => \N__21690\
        );

    \I__1961\ : InMux
    port map (
            O => \N__21690\,
            I => \N__21687\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__21687\,
            I => \N__21684\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__21684\,
            I => \N__21681\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__21681\,
            I => \current_shift_inst.PI_CTRL.integrator_1_22\
        );

    \I__1957\ : InMux
    port map (
            O => \N__21678\,
            I => \N__21675\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__21675\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__1955\ : InMux
    port map (
            O => \N__21672\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__21669\,
            I => \N__21666\
        );

    \I__1953\ : InMux
    port map (
            O => \N__21666\,
            I => \N__21663\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__21663\,
            I => \N__21660\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__21660\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__1950\ : InMux
    port map (
            O => \N__21657\,
            I => \N__21654\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__21654\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__1948\ : InMux
    port map (
            O => \N__21651\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__21648\,
            I => \N__21645\
        );

    \I__1946\ : InMux
    port map (
            O => \N__21645\,
            I => \N__21642\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__21642\,
            I => \N__21639\
        );

    \I__1944\ : Span4Mux_h
    port map (
            O => \N__21639\,
            I => \N__21636\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__21636\,
            I => \current_shift_inst.PI_CTRL.integrator_1_8\
        );

    \I__1942\ : InMux
    port map (
            O => \N__21633\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__21630\,
            I => \N__21627\
        );

    \I__1940\ : InMux
    port map (
            O => \N__21627\,
            I => \N__21624\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__21624\,
            I => \N__21621\
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__21621\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__1937\ : InMux
    port map (
            O => \N__21618\,
            I => \N__21615\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__21615\,
            I => \N__21612\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__21612\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__1934\ : InMux
    port map (
            O => \N__21609\,
            I => \bfn_2_11_0_\
        );

    \I__1933\ : InMux
    port map (
            O => \N__21606\,
            I => \N__21603\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__21603\,
            I => \N__21600\
        );

    \I__1931\ : Odrv12
    port map (
            O => \N__21600\,
            I => \current_shift_inst.PI_CTRL.integrator_1_10\
        );

    \I__1930\ : InMux
    port map (
            O => \N__21597\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__21594\,
            I => \N__21591\
        );

    \I__1928\ : InMux
    port map (
            O => \N__21591\,
            I => \N__21588\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__21588\,
            I => \N__21585\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__21585\,
            I => \current_shift_inst.PI_CTRL.integrator_1_11\
        );

    \I__1925\ : InMux
    port map (
            O => \N__21582\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__1924\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21576\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__21576\,
            I => \N__21573\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__21573\,
            I => \current_shift_inst.PI_CTRL.integrator_1_12\
        );

    \I__1921\ : InMux
    port map (
            O => \N__21570\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__21567\,
            I => \N__21564\
        );

    \I__1919\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21561\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__21561\,
            I => \N__21558\
        );

    \I__1917\ : Odrv12
    port map (
            O => \N__21558\,
            I => \current_shift_inst.PI_CTRL.integrator_1_13\
        );

    \I__1916\ : InMux
    port map (
            O => \N__21555\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__21552\,
            I => \N__21549\
        );

    \I__1914\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21546\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__21546\,
            I => \N__21543\
        );

    \I__1912\ : Odrv12
    port map (
            O => \N__21543\,
            I => \current_shift_inst.PI_CTRL.integrator_1_14\
        );

    \I__1911\ : InMux
    port map (
            O => \N__21540\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__1910\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21534\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__21534\,
            I => \N__21531\
        );

    \I__1908\ : Span4Mux_h
    port map (
            O => \N__21531\,
            I => \N__21528\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__21528\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_15\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__21525\,
            I => \N__21519\
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__21524\,
            I => \N__21515\
        );

    \I__1904\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21512\
        );

    \I__1903\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21496\
        );

    \I__1902\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21496\
        );

    \I__1901\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21496\
        );

    \I__1900\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21496\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__21512\,
            I => \N__21493\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__21511\,
            I => \N__21490\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__21510\,
            I => \N__21487\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__21509\,
            I => \N__21484\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__21508\,
            I => \N__21481\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__21507\,
            I => \N__21478\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__21506\,
            I => \N__21475\
        );

    \I__1892\ : CascadeMux
    port map (
            O => \N__21505\,
            I => \N__21472\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__21496\,
            I => \N__21469\
        );

    \I__1890\ : Span4Mux_h
    port map (
            O => \N__21493\,
            I => \N__21466\
        );

    \I__1889\ : InMux
    port map (
            O => \N__21490\,
            I => \N__21459\
        );

    \I__1888\ : InMux
    port map (
            O => \N__21487\,
            I => \N__21459\
        );

    \I__1887\ : InMux
    port map (
            O => \N__21484\,
            I => \N__21459\
        );

    \I__1886\ : InMux
    port map (
            O => \N__21481\,
            I => \N__21450\
        );

    \I__1885\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21450\
        );

    \I__1884\ : InMux
    port map (
            O => \N__21475\,
            I => \N__21450\
        );

    \I__1883\ : InMux
    port map (
            O => \N__21472\,
            I => \N__21450\
        );

    \I__1882\ : Span4Mux_v
    port map (
            O => \N__21469\,
            I => \N__21447\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__21466\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__21459\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__21450\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__21447\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__21438\,
            I => \N__21435\
        );

    \I__1876\ : InMux
    port map (
            O => \N__21435\,
            I => \N__21432\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__21432\,
            I => \N__21429\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__21429\,
            I => \current_shift_inst.PI_CTRL.un1_integrator\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__21426\,
            I => \N__21423\
        );

    \I__1872\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21420\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__21420\,
            I => \N__21417\
        );

    \I__1870\ : Odrv12
    port map (
            O => \N__21417\,
            I => \current_shift_inst.PI_CTRL.integrator_1_2\
        );

    \I__1869\ : InMux
    port map (
            O => \N__21414\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__21411\,
            I => \N__21408\
        );

    \I__1867\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21405\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__21405\,
            I => \N__21402\
        );

    \I__1865\ : Odrv12
    port map (
            O => \N__21402\,
            I => \current_shift_inst.PI_CTRL.integrator_1_3\
        );

    \I__1864\ : InMux
    port map (
            O => \N__21399\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__21396\,
            I => \N__21393\
        );

    \I__1862\ : InMux
    port map (
            O => \N__21393\,
            I => \N__21390\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__21390\,
            I => \N__21387\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__21387\,
            I => \current_shift_inst.PI_CTRL.integrator_1_4\
        );

    \I__1859\ : InMux
    port map (
            O => \N__21384\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__21381\,
            I => \N__21378\
        );

    \I__1857\ : InMux
    port map (
            O => \N__21378\,
            I => \N__21375\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__21375\,
            I => \N__21372\
        );

    \I__1855\ : Odrv12
    port map (
            O => \N__21372\,
            I => \current_shift_inst.PI_CTRL.integrator_1_5\
        );

    \I__1854\ : InMux
    port map (
            O => \N__21369\,
            I => \N__21366\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__21366\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__1852\ : InMux
    port map (
            O => \N__21363\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__21360\,
            I => \N__21357\
        );

    \I__1850\ : InMux
    port map (
            O => \N__21357\,
            I => \N__21354\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__21354\,
            I => \N__21351\
        );

    \I__1848\ : Span4Mux_h
    port map (
            O => \N__21351\,
            I => \N__21348\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__21348\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__1846\ : InMux
    port map (
            O => \N__21345\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__1845\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21339\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__21339\,
            I => \N__21336\
        );

    \I__1843\ : Span4Mux_v
    port map (
            O => \N__21336\,
            I => \N__21333\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__21333\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_14\
        );

    \I__1841\ : InMux
    port map (
            O => \N__21330\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\
        );

    \I__1840\ : InMux
    port map (
            O => \N__21327\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\
        );

    \I__1839\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21321\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__21321\,
            I => \N_94_i_i\
        );

    \I__1837\ : InMux
    port map (
            O => \N__21318\,
            I => \N__21315\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__21315\,
            I => \N__21312\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__21312\,
            I => \N__21309\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__21309\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_6\
        );

    \I__1833\ : InMux
    port map (
            O => \N__21306\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__21303\,
            I => \N__21300\
        );

    \I__1831\ : InMux
    port map (
            O => \N__21300\,
            I => \N__21297\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__21297\,
            I => \N__21294\
        );

    \I__1829\ : Span4Mux_v
    port map (
            O => \N__21294\,
            I => \N__21291\
        );

    \I__1828\ : Odrv4
    port map (
            O => \N__21291\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_7\
        );

    \I__1827\ : InMux
    port map (
            O => \N__21288\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\
        );

    \I__1826\ : InMux
    port map (
            O => \N__21285\,
            I => \N__21282\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__21282\,
            I => \N__21279\
        );

    \I__1824\ : Span4Mux_v
    port map (
            O => \N__21279\,
            I => \N__21276\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__21276\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_8\
        );

    \I__1822\ : InMux
    port map (
            O => \N__21273\,
            I => \bfn_1_11_0_\
        );

    \I__1821\ : InMux
    port map (
            O => \N__21270\,
            I => \N__21267\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__21267\,
            I => \N__21264\
        );

    \I__1819\ : Span4Mux_v
    port map (
            O => \N__21264\,
            I => \N__21261\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__21261\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_9\
        );

    \I__1817\ : InMux
    port map (
            O => \N__21258\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\
        );

    \I__1816\ : InMux
    port map (
            O => \N__21255\,
            I => \N__21252\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__21252\,
            I => \N__21249\
        );

    \I__1814\ : Span4Mux_v
    port map (
            O => \N__21249\,
            I => \N__21246\
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__21246\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_10\
        );

    \I__1812\ : InMux
    port map (
            O => \N__21243\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\
        );

    \I__1811\ : InMux
    port map (
            O => \N__21240\,
            I => \N__21237\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__21237\,
            I => \N__21234\
        );

    \I__1809\ : Span4Mux_v
    port map (
            O => \N__21234\,
            I => \N__21231\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__21231\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_11\
        );

    \I__1807\ : InMux
    port map (
            O => \N__21228\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\
        );

    \I__1806\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21222\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__21222\,
            I => \N__21219\
        );

    \I__1804\ : Span4Mux_v
    port map (
            O => \N__21219\,
            I => \N__21216\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__21216\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_12\
        );

    \I__1802\ : InMux
    port map (
            O => \N__21213\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\
        );

    \I__1801\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21207\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__21207\,
            I => \N__21204\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__21204\,
            I => \N__21201\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__21201\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_13\
        );

    \I__1797\ : InMux
    port map (
            O => \N__21198\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\
        );

    \I__1796\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21192\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__21192\,
            I => \N__21189\
        );

    \I__1794\ : Span4Mux_v
    port map (
            O => \N__21189\,
            I => \N__21186\
        );

    \I__1793\ : Odrv4
    port map (
            O => \N__21186\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_0\
        );

    \I__1792\ : CascadeMux
    port map (
            O => \N__21183\,
            I => \N__21180\
        );

    \I__1791\ : InMux
    port map (
            O => \N__21180\,
            I => \N__21177\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__21177\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_15\
        );

    \I__1789\ : InMux
    port map (
            O => \N__21174\,
            I => \N__21171\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__21171\,
            I => \N__21168\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__21168\,
            I => \N__21165\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__21165\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_1\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__21162\,
            I => \N__21159\
        );

    \I__1784\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21156\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__21156\,
            I => \N__21153\
        );

    \I__1782\ : Odrv4
    port map (
            O => \N__21153\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_16\
        );

    \I__1781\ : InMux
    port map (
            O => \N__21150\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\
        );

    \I__1780\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21144\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__21144\,
            I => \N__21141\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__21141\,
            I => \N__21138\
        );

    \I__1777\ : Odrv4
    port map (
            O => \N__21138\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_2\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__21135\,
            I => \N__21132\
        );

    \I__1775\ : InMux
    port map (
            O => \N__21132\,
            I => \N__21129\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__21129\,
            I => \N__21126\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__21126\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_17\
        );

    \I__1772\ : InMux
    port map (
            O => \N__21123\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\
        );

    \I__1771\ : InMux
    port map (
            O => \N__21120\,
            I => \N__21117\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__21117\,
            I => \N__21114\
        );

    \I__1769\ : Span4Mux_v
    port map (
            O => \N__21114\,
            I => \N__21111\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__21111\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_3\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__21108\,
            I => \N__21105\
        );

    \I__1766\ : InMux
    port map (
            O => \N__21105\,
            I => \N__21102\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__21102\,
            I => \N__21099\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__21099\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_18\
        );

    \I__1763\ : InMux
    port map (
            O => \N__21096\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\
        );

    \I__1762\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21090\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__21090\,
            I => \N__21087\
        );

    \I__1760\ : Span4Mux_v
    port map (
            O => \N__21087\,
            I => \N__21084\
        );

    \I__1759\ : Odrv4
    port map (
            O => \N__21084\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_4\
        );

    \I__1758\ : InMux
    port map (
            O => \N__21081\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__21078\,
            I => \N__21075\
        );

    \I__1756\ : InMux
    port map (
            O => \N__21075\,
            I => \N__21072\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__21072\,
            I => \N__21069\
        );

    \I__1754\ : Span4Mux_v
    port map (
            O => \N__21069\,
            I => \N__21066\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__21066\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_5\
        );

    \I__1752\ : InMux
    port map (
            O => \N__21063\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\
        );

    \I__1751\ : IoInMux
    port map (
            O => \N__21060\,
            I => \N__21057\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__21057\,
            I => \N__21054\
        );

    \I__1749\ : Span4Mux_s3_v
    port map (
            O => \N__21054\,
            I => \N__21051\
        );

    \I__1748\ : Span4Mux_h
    port map (
            O => \N__21051\,
            I => \N__21048\
        );

    \I__1747\ : Sp12to4
    port map (
            O => \N__21048\,
            I => \N__21045\
        );

    \I__1746\ : Span12Mux_v
    port map (
            O => \N__21045\,
            I => \N__21042\
        );

    \I__1745\ : Span12Mux_v
    port map (
            O => \N__21042\,
            I => \N__21039\
        );

    \I__1744\ : Odrv12
    port map (
            O => \N__21039\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1743\ : IoInMux
    port map (
            O => \N__21036\,
            I => \N__21033\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__21033\,
            I => \N__21030\
        );

    \I__1741\ : IoSpan4Mux
    port map (
            O => \N__21030\,
            I => \N__21027\
        );

    \I__1740\ : IoSpan4Mux
    port map (
            O => \N__21027\,
            I => \N__21024\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__21024\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_15_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_28_0_\
        );

    \IN_MUX_bfv_15_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_15_29_0_\
        );

    \IN_MUX_bfv_15_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_15_30_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_8_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_8_22_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_11_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryinitout => \bfn_11_21_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_16_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_28_0_\
        );

    \IN_MUX_bfv_16_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_16_29_0_\
        );

    \IN_MUX_bfv_16_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            carryinitout => \bfn_16_30_0_\
        );

    \IN_MUX_bfv_17_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_26_0_\
        );

    \IN_MUX_bfv_17_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_0_cry_7\,
            carryinitout => \bfn_17_27_0_\
        );

    \IN_MUX_bfv_20_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_25_0_\
        );

    \IN_MUX_bfv_20_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_7\,
            carryinitout => \bfn_20_26_0_\
        );

    \IN_MUX_bfv_20_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_15\,
            carryinitout => \bfn_20_27_0_\
        );

    \IN_MUX_bfv_17_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_24_0_\
        );

    \IN_MUX_bfv_17_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_17_25_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_16_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_16_24_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_7\,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_15\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_30\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_10_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_7_0_\
        );

    \IN_MUX_bfv_10_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.counter_cry_7\,
            carryinitout => \bfn_10_8_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.counter_cry_15\,
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.counter_cry_23\,
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_7\,
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_15\,
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_30\,
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.counter_cry_7\,
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.counter_cry_15\,
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.counter_cry_23\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_11_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_25_0_\
        );

    \IN_MUX_bfv_11_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_7\,
            carryinitout => \bfn_11_26_0_\
        );

    \IN_MUX_bfv_11_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_15\,
            carryinitout => \bfn_11_27_0_\
        );

    \IN_MUX_bfv_11_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_30\,
            carryinitout => \bfn_11_28_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8\,
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16\,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24\,
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7\,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_13_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15\,
            carryinitout => \bfn_13_21_0_\
        );

    \IN_MUX_bfv_13_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23\,
            carryinitout => \bfn_13_22_0_\
        );

    \IN_MUX_bfv_12_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_27_0_\
        );

    \IN_MUX_bfv_12_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.counter_cry_7\,
            carryinitout => \bfn_12_28_0_\
        );

    \IN_MUX_bfv_12_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.counter_cry_15\,
            carryinitout => \bfn_12_29_0_\
        );

    \IN_MUX_bfv_12_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.counter_cry_23\,
            carryinitout => \bfn_12_30_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_7\,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_15\,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_30\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16\,
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24\,
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7\,
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15\,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.counter_cry_7\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.counter_cry_15\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.counter_cry_23\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_14_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_14_25_0_\
        );

    \IN_MUX_bfv_14_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_14_26_0_\
        );

    \IN_MUX_bfv_14_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_14_27_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_13_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_13_25_0_\
        );

    \IN_MUX_bfv_13_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_13_26_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_17_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_17_21_0_\
        );

    \IN_MUX_bfv_17_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_17_22_0_\
        );

    \IN_MUX_bfv_17_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_17_23_0_\
        );

    \IN_MUX_bfv_3_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_11_0_\
        );

    \IN_MUX_bfv_3_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_3_12_0_\
        );

    \IN_MUX_bfv_3_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_15\,
            carryinitout => \bfn_3_13_0_\
        );

    \IN_MUX_bfv_3_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_23\,
            carryinitout => \bfn_3_14_0_\
        );

    \IN_MUX_bfv_10_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_20_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_10_23_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            carryinitout => \bfn_5_14_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21060\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21036\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__31470\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst1.stoper_tr.un2_start_0_g\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__28083\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_tr.un2_start_0_g\
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__38226\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_153_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__46576\,
            CLKHFEN => \N__46578\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__46577\,
            RGB2PWM => \N__21324\,
            RGB1 => rgb_g_wire,
            CURREN => \N__46828\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__22140\,
            RGB0PWM => \N__52089\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__31641\,
            in1 => \N__21369\,
            in2 => \_gnd_net_\,
            in3 => \N__22597\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52500\,
            ce => 'H',
            sr => \N__51989\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__22596\,
            in1 => \N__21618\,
            in2 => \_gnd_net_\,
            in3 => \N__31642\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52500\,
            ce => 'H',
            sr => \N__51989\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21195\,
            in2 => \N__21183\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_16\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21174\,
            in2 => \N__21162\,
            in3 => \N__21150\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21147\,
            in2 => \N__21135\,
            in3 => \N__21123\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21120\,
            in2 => \N__21108\,
            in3 => \N__21096\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21093\,
            in2 => \N__21524\,
            in3 => \N__21081\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21518\,
            in2 => \N__21078\,
            in3 => \N__21063\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21318\,
            in2 => \N__21525\,
            in3 => \N__21306\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21522\,
            in2 => \N__21303\,
            in3 => \N__21288\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21285\,
            in2 => \N__21505\,
            in3 => \N__21273\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_24\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21270\,
            in2 => \N__21509\,
            in3 => \N__21258\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21255\,
            in2 => \N__21506\,
            in3 => \N__21243\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21240\,
            in2 => \N__21510\,
            in3 => \N__21228\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21225\,
            in2 => \N__21507\,
            in3 => \N__21213\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21210\,
            in2 => \N__21511\,
            in3 => \N__21198\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21342\,
            in2 => \N__21508\,
            in3 => \N__21330\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21327\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22621\,
            in1 => \N__31589\,
            in2 => \_gnd_net_\,
            in3 => \N__21768\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52494\,
            ce => 'H',
            sr => \N__52007\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22622\,
            in1 => \N__31590\,
            in2 => \_gnd_net_\,
            in3 => \N__21678\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52494\,
            ce => 'H',
            sr => \N__52007\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31588\,
            in1 => \N__22623\,
            in2 => \_gnd_net_\,
            in3 => \N__21954\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52494\,
            ce => 'H',
            sr => \N__52007\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22624\,
            in1 => \N__31592\,
            in2 => \_gnd_net_\,
            in3 => \N__21702\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52491\,
            ce => 'H',
            sr => \N__52014\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22625\,
            in1 => \N__31593\,
            in2 => \_gnd_net_\,
            in3 => \N__21933\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52491\,
            ce => 'H',
            sr => \N__52014\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22626\,
            in1 => \N__31594\,
            in2 => \_gnd_net_\,
            in3 => \N__21873\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52491\,
            ce => 'H',
            sr => \N__52014\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31591\,
            in1 => \N__22646\,
            in2 => \_gnd_net_\,
            in3 => \N__21840\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52485\,
            ce => 'H',
            sr => \N__52023\
        );

    \phase_controller_inst1.N_94_i_i_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__52088\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36612\,
            lcout => \N_94_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21537\,
            in2 => \_gnd_net_\,
            in3 => \N__21523\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30232\,
            in1 => \N__30106\,
            in2 => \N__30928\,
            in3 => \N__30173\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__31643\,
            in1 => \N__21657\,
            in2 => \_gnd_net_\,
            in3 => \N__22595\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52499\,
            ce => 'H',
            sr => \N__51980\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36681\,
            in2 => \N__21438\,
            in3 => \N__22628\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \N__52497\,
            ce => 'H',
            sr => \N__51991\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__22627\,
            in1 => \N__30427\,
            in2 => \N__21426\,
            in3 => \N__21414\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \N__52497\,
            ce => 'H',
            sr => \N__51991\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__22647\,
            in1 => \N__30351\,
            in2 => \N__21411\,
            in3 => \N__21399\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \N__52497\,
            ce => 'H',
            sr => \N__51991\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30295\,
            in2 => \N__21396\,
            in3 => \N__21384\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30228\,
            in2 => \N__21381\,
            in3 => \N__21363\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30171\,
            in2 => \N__21360\,
            in3 => \N__21345\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30105\,
            in2 => \N__21669\,
            in3 => \N__21651\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30057\,
            in2 => \N__21648\,
            in3 => \N__21633\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30927\,
            in2 => \N__21630\,
            in3 => \N__21609\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21606\,
            in2 => \N__30860\,
            in3 => \N__21597\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30793\,
            in2 => \N__21594\,
            in3 => \N__21582\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21579\,
            in2 => \N__30731\,
            in3 => \N__21570\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30655\,
            in2 => \N__21567\,
            in3 => \N__21555\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30598\,
            in2 => \N__21552\,
            in3 => \N__21540\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30547\,
            in2 => \N__21813\,
            in3 => \N__21798\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30478\,
            in2 => \N__21795\,
            in3 => \N__21786\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31419\,
            in2 => \N__21783\,
            in3 => \N__21762\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31360\,
            in2 => \N__21759\,
            in3 => \N__21747\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31296\,
            in2 => \N__21744\,
            in3 => \N__21729\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21726\,
            in2 => \N__31229\,
            in3 => \N__21717\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31155\,
            in2 => \N__21714\,
            in3 => \N__21696\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31101\,
            in2 => \N__21693\,
            in3 => \N__21672\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31041\,
            in2 => \N__21966\,
            in3 => \N__21948\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30981\,
            in2 => \N__21945\,
            in3 => \N__21927\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32016\,
            in2 => \N__21924\,
            in3 => \N__21909\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31954\,
            in2 => \N__21906\,
            in3 => \N__21891\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31878\,
            in2 => \N__21888\,
            in3 => \N__21867\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21864\,
            in2 => \N__31824\,
            in3 => \N__21855\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31747\,
            in2 => \N__21852\,
            in3 => \N__21834\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31689\,
            in2 => \N__21831\,
            in3 => \N__21816\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_er_31_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22077\,
            in1 => \N__31595\,
            in2 => \N__22068\,
            in3 => \N__22053\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52486\,
            ce => \N__22649\,
            sr => \N__52008\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31582\,
            in1 => \N__22632\,
            in2 => \_gnd_net_\,
            in3 => \N__22050\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52482\,
            ce => 'H',
            sr => \N__52015\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__22041\,
            in1 => \N__31587\,
            in2 => \N__22652\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52482\,
            ce => 'H',
            sr => \N__52015\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__22032\,
            in1 => \_gnd_net_\,
            in2 => \N__22653\,
            in3 => \N__31584\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52482\,
            ce => 'H',
            sr => \N__52015\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31583\,
            in1 => \N__22633\,
            in2 => \_gnd_net_\,
            in3 => \N__22023\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52482\,
            ce => 'H',
            sr => \N__52015\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__22017\,
            in1 => \N__31586\,
            in2 => \N__22651\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52482\,
            ce => 'H',
            sr => \N__52015\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__22011\,
            in1 => \N__31585\,
            in2 => \N__22650\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52482\,
            ce => 'H',
            sr => \N__52015\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31613\,
            in1 => \N__22002\,
            in2 => \_gnd_net_\,
            in3 => \N__22648\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52478\,
            ce => 'H',
            sr => \N__52024\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21993\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.un8_start_stop_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__52087\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36611\,
            lcout => un8_start_stop,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22550\,
            in1 => \N__31650\,
            in2 => \_gnd_net_\,
            in3 => \N__22131\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52498\,
            ce => 'H',
            sr => \N__51976\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__31648\,
            in1 => \_gnd_net_\,
            in2 => \N__22122\,
            in3 => \N__22552\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52498\,
            ce => 'H',
            sr => \N__51976\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31647\,
            in1 => \N__22113\,
            in2 => \_gnd_net_\,
            in3 => \N__22551\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52498\,
            ce => 'H',
            sr => \N__51976\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__31649\,
            in1 => \N__22104\,
            in2 => \_gnd_net_\,
            in3 => \N__22553\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52498\,
            ce => 'H',
            sr => \N__51976\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22554\,
            in1 => \N__31652\,
            in2 => \_gnd_net_\,
            in3 => \N__22098\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52495\,
            ce => 'H',
            sr => \N__51981\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31651\,
            in1 => \N__22092\,
            in2 => \_gnd_net_\,
            in3 => \N__22557\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52495\,
            ce => 'H',
            sr => \N__51981\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22555\,
            in1 => \N__31653\,
            in2 => \_gnd_net_\,
            in3 => \N__22086\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52495\,
            ce => 'H',
            sr => \N__51981\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22244\,
            in2 => \_gnd_net_\,
            in3 => \N__23673\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52495\,
            ce => 'H',
            sr => \N__51981\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__22556\,
            in1 => \N__31654\,
            in2 => \_gnd_net_\,
            in3 => \N__22170\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52495\,
            ce => 'H',
            sr => \N__51981\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23669\,
            in2 => \N__22245\,
            in3 => \N__22243\,
            lcout => \current_shift_inst.control_input_1\,
            ltout => OPEN,
            carryin => \bfn_3_11_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23688\,
            in2 => \_gnd_net_\,
            in3 => \N__22164\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22359\,
            in2 => \_gnd_net_\,
            in3 => \N__22161\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23649\,
            in2 => \_gnd_net_\,
            in3 => \N__22158\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23634\,
            in2 => \_gnd_net_\,
            in3 => \N__22155\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22365\,
            in2 => \_gnd_net_\,
            in3 => \N__22152\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22395\,
            in2 => \_gnd_net_\,
            in3 => \N__22149\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22371\,
            in2 => \_gnd_net_\,
            in3 => \N__22146\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22377\,
            in2 => \_gnd_net_\,
            in3 => \N__22143\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_12_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23586\,
            in2 => \_gnd_net_\,
            in3 => \N__22197\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22455\,
            in2 => \_gnd_net_\,
            in3 => \N__22194\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23598\,
            in2 => \_gnd_net_\,
            in3 => \N__22191\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22353\,
            in2 => \_gnd_net_\,
            in3 => \N__22188\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22449\,
            in2 => \_gnd_net_\,
            in3 => \N__22185\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_12\,
            carryout => \current_shift_inst.control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23574\,
            in2 => \_gnd_net_\,
            in3 => \N__22182\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_13\,
            carryout => \current_shift_inst.control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23529\,
            in2 => \_gnd_net_\,
            in3 => \N__22179\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_14\,
            carryout => \current_shift_inst.control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23700\,
            in2 => \_gnd_net_\,
            in3 => \N__22176\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_3_13_0_\,
            carryout => \current_shift_inst.control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23541\,
            in2 => \_gnd_net_\,
            in3 => \N__22173\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_16\,
            carryout => \current_shift_inst.control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22443\,
            in2 => \_gnd_net_\,
            in3 => \N__22224\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_17\,
            carryout => \current_shift_inst.control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23931\,
            in2 => \_gnd_net_\,
            in3 => \N__22221\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_18\,
            carryout => \current_shift_inst.control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22437\,
            in2 => \_gnd_net_\,
            in3 => \N__22218\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_19\,
            carryout => \current_shift_inst.control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23553\,
            in2 => \_gnd_net_\,
            in3 => \N__22215\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_20\,
            carryout => \current_shift_inst.control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22407\,
            in2 => \_gnd_net_\,
            in3 => \N__22212\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_21\,
            carryout => \current_shift_inst.control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22719\,
            in2 => \_gnd_net_\,
            in3 => \N__22209\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_22\,
            carryout => \current_shift_inst.control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22401\,
            in2 => \_gnd_net_\,
            in3 => \N__22206\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_3_14_0_\,
            carryout => \current_shift_inst.control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22713\,
            in2 => \_gnd_net_\,
            in3 => \N__22203\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_24\,
            carryout => \current_shift_inst.control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23562\,
            in2 => \_gnd_net_\,
            in3 => \N__22200\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_25\,
            carryout => \current_shift_inst.control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22413\,
            in2 => \_gnd_net_\,
            in3 => \N__22284\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_26\,
            carryout => \current_shift_inst.control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24414\,
            in2 => \_gnd_net_\,
            in3 => \N__22281\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_27\,
            carryout => \current_shift_inst.control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22695\,
            in2 => \_gnd_net_\,
            in3 => \N__22278\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_28\,
            carryout => \current_shift_inst.control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__24586\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22275\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => \current_shift_inst.control_input_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22272\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31635\,
            in1 => \N__22269\,
            in2 => \_gnd_net_\,
            in3 => \N__22620\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52470\,
            ce => 'H',
            sr => \N__52016\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__30059\,
            in1 => \N__30296\,
            in2 => \N__30368\,
            in3 => \N__22257\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__22686\,
            in1 => \N__22299\,
            in2 => \N__22248\,
            in3 => \N__22314\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24560\,
            lcout => \current_shift_inst.N_1571_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30597\,
            in1 => \N__30651\,
            in2 => \N__30794\,
            in3 => \N__30462\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__30113\,
            in1 => \N__30172\,
            in2 => \_gnd_net_\,
            in3 => \N__30239\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__30058\,
            in1 => \N__30929\,
            in2 => \N__22335\,
            in3 => \N__22332\,
            lcout => \current_shift_inst.PI_CTRL.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010111"
        )
    port map (
            in0 => \N__30352\,
            in1 => \N__30431\,
            in2 => \N__36697\,
            in3 => \N__30294\,
            lcout => \current_shift_inst.PI_CTRL.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__30853\,
            in1 => \N__22389\,
            in2 => \N__30548\,
            in3 => \N__22290\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__31636\,
            in1 => \N__31350\,
            in2 => \N__22326\,
            in3 => \N__22461\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22707\,
            in1 => \N__22422\,
            in2 => \N__22323\,
            in3 => \N__22320\,
            lcout => \current_shift_inst.PI_CTRL.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22431\,
            in1 => \N__22383\,
            in2 => \N__22347\,
            in3 => \N__22305\,
            lcout => \current_shift_inst.PI_CTRL.N_46_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31227\,
            in1 => \N__31429\,
            in2 => \N__31307\,
            in3 => \N__31114\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__24639\,
            in1 => \N__24135\,
            in2 => \_gnd_net_\,
            in3 => \N__24563\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31756\,
            in2 => \_gnd_net_\,
            in3 => \N__31042\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31757\,
            in1 => \N__30540\,
            in2 => \N__31049\,
            in3 => \N__30852\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__24565\,
            in1 => \N__24858\,
            in2 => \_gnd_net_\,
            in3 => \N__24111\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__24615\,
            in1 => \N__24123\,
            in2 => \_gnd_net_\,
            in3 => \N__24564\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__24562\,
            in1 => \N__24147\,
            in2 => \_gnd_net_\,
            in3 => \N__24654\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__24003\,
            in1 => \N__24693\,
            in2 => \_gnd_net_\,
            in3 => \N__24561\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110101"
        )
    port map (
            in0 => \N__24792\,
            in1 => \_gnd_net_\,
            in2 => \N__24587\,
            in3 => \N__24267\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31825\,
            in1 => \N__31882\,
            in2 => \N__31706\,
            in3 => \N__30727\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100011011"
        )
    port map (
            in0 => \N__24588\,
            in1 => \N__24825\,
            in2 => \N__24090\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100110101"
        )
    port map (
            in0 => \N__24774\,
            in1 => \N__24252\,
            in2 => \N__24594\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__24592\,
            in1 => \N__24192\,
            in2 => \_gnd_net_\,
            in3 => \N__24996\,
            lcout => \current_shift_inst.control_input_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__24963\,
            in1 => \N__24381\,
            in2 => \_gnd_net_\,
            in3 => \N__24593\,
            lcout => \current_shift_inst.control_input_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31156\,
            in1 => \N__32017\,
            in2 => \N__31958\,
            in3 => \N__30982\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32018\,
            in1 => \N__31953\,
            in2 => \N__30989\,
            in3 => \N__31157\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__24288\,
            in1 => \N__24585\,
            in2 => \_gnd_net_\,
            in3 => \N__25098\,
            lcout => \current_shift_inst.control_input_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__24348\,
            in1 => \N__24921\,
            in2 => \_gnd_net_\,
            in3 => \N__24581\,
            lcout => \current_shift_inst.control_input_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__24583\,
            in1 => \N__24882\,
            in2 => \_gnd_net_\,
            in3 => \N__24324\,
            lcout => \current_shift_inst.control_input_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__24582\,
            in1 => \N__24336\,
            in2 => \_gnd_net_\,
            in3 => \N__24903\,
            lcout => \current_shift_inst.control_input_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__25146\,
            in1 => \N__24309\,
            in2 => \_gnd_net_\,
            in3 => \N__24584\,
            lcout => \current_shift_inst.control_input_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31690\,
            in1 => \N__31886\,
            in2 => \N__31826\,
            in3 => \N__30723\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24559\,
            lcout => \current_shift_inst.control_input_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31228\,
            in1 => \N__31303\,
            in2 => \N__31436\,
            in3 => \N__31115\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_46_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31640\,
            in2 => \N__22689\,
            in3 => \N__31361\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22677\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52449\,
            ce => 'H',
            sr => \N__52031\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31655\,
            in1 => \N__22558\,
            in2 => \_gnd_net_\,
            in3 => \N__22473\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52492\,
            ce => 'H',
            sr => \N__51970\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30602\,
            in1 => \N__30656\,
            in2 => \N__30482\,
            in3 => \N__30774\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22824\,
            in2 => \_gnd_net_\,
            in3 => \N__22833\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22818\,
            in2 => \_gnd_net_\,
            in3 => \N__22809\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__52483\,
            ce => 'H',
            sr => \N__51977\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22806\,
            in3 => \N__22794\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__52483\,
            ce => 'H',
            sr => \N__51977\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22791\,
            in2 => \_gnd_net_\,
            in3 => \N__22782\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__52483\,
            ce => 'H',
            sr => \N__51977\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22779\,
            in2 => \_gnd_net_\,
            in3 => \N__22770\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__52483\,
            ce => 'H',
            sr => \N__51977\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22767\,
            in2 => \_gnd_net_\,
            in3 => \N__22758\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__52483\,
            ce => 'H',
            sr => \N__51977\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22755\,
            in2 => \_gnd_net_\,
            in3 => \N__22746\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__52483\,
            ce => 'H',
            sr => \N__51977\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22743\,
            in2 => \_gnd_net_\,
            in3 => \N__22734\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__52483\,
            ce => 'H',
            sr => \N__51977\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22731\,
            in2 => \_gnd_net_\,
            in3 => \N__22722\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__52479\,
            ce => 'H',
            sr => \N__51982\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22932\,
            in2 => \_gnd_net_\,
            in3 => \N__22923\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__52479\,
            ce => 'H',
            sr => \N__51982\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22920\,
            in2 => \_gnd_net_\,
            in3 => \N__22911\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__52479\,
            ce => 'H',
            sr => \N__51982\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22908\,
            in3 => \N__22896\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__52479\,
            ce => 'H',
            sr => \N__51982\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22893\,
            in2 => \_gnd_net_\,
            in3 => \N__22884\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__52479\,
            ce => 'H',
            sr => \N__51982\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22881\,
            in2 => \_gnd_net_\,
            in3 => \N__22872\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__52479\,
            ce => 'H',
            sr => \N__51982\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22869\,
            in2 => \_gnd_net_\,
            in3 => \N__22860\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            clk => \N__52479\,
            ce => 'H',
            sr => \N__51982\
        );

    \current_shift_inst.PI_CTRL.error_control_15_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22857\,
            in2 => \_gnd_net_\,
            in3 => \N__22848\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            clk => \N__52479\,
            ce => 'H',
            sr => \N__51982\
        );

    \current_shift_inst.PI_CTRL.error_control_16_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22845\,
            in2 => \_gnd_net_\,
            in3 => \N__22836\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_16\,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            clk => \N__52471\,
            ce => 'H',
            sr => \N__51992\
        );

    \current_shift_inst.PI_CTRL.error_control_17_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23040\,
            in2 => \_gnd_net_\,
            in3 => \N__23031\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            clk => \N__52471\,
            ce => 'H',
            sr => \N__51992\
        );

    \current_shift_inst.PI_CTRL.error_control_18_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23028\,
            in2 => \_gnd_net_\,
            in3 => \N__23019\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            clk => \N__52471\,
            ce => 'H',
            sr => \N__51992\
        );

    \current_shift_inst.PI_CTRL.error_control_19_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23016\,
            in2 => \_gnd_net_\,
            in3 => \N__23007\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            clk => \N__52471\,
            ce => 'H',
            sr => \N__51992\
        );

    \current_shift_inst.PI_CTRL.error_control_20_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23004\,
            in2 => \_gnd_net_\,
            in3 => \N__22995\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            clk => \N__52471\,
            ce => 'H',
            sr => \N__51992\
        );

    \current_shift_inst.PI_CTRL.error_control_21_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22992\,
            in2 => \_gnd_net_\,
            in3 => \N__22983\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            clk => \N__52471\,
            ce => 'H',
            sr => \N__51992\
        );

    \current_shift_inst.PI_CTRL.error_control_22_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22980\,
            in2 => \_gnd_net_\,
            in3 => \N__22971\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            clk => \N__52471\,
            ce => 'H',
            sr => \N__51992\
        );

    \current_shift_inst.PI_CTRL.error_control_23_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22968\,
            in3 => \N__22956\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            clk => \N__52471\,
            ce => 'H',
            sr => \N__51992\
        );

    \current_shift_inst.PI_CTRL.error_control_24_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22953\,
            in2 => \_gnd_net_\,
            in3 => \N__22944\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_24\,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            clk => \N__52465\,
            ce => 'H',
            sr => \N__51995\
        );

    \current_shift_inst.PI_CTRL.error_control_25_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22941\,
            in2 => \_gnd_net_\,
            in3 => \N__23163\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            clk => \N__52465\,
            ce => 'H',
            sr => \N__51995\
        );

    \current_shift_inst.PI_CTRL.error_control_26_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23160\,
            in2 => \_gnd_net_\,
            in3 => \N__23151\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            clk => \N__52465\,
            ce => 'H',
            sr => \N__51995\
        );

    \current_shift_inst.PI_CTRL.error_control_27_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23148\,
            in2 => \_gnd_net_\,
            in3 => \N__23139\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            clk => \N__52465\,
            ce => 'H',
            sr => \N__51995\
        );

    \current_shift_inst.PI_CTRL.error_control_28_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23136\,
            in2 => \_gnd_net_\,
            in3 => \N__23127\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            clk => \N__52465\,
            ce => 'H',
            sr => \N__51995\
        );

    \current_shift_inst.PI_CTRL.error_control_29_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23124\,
            in2 => \_gnd_net_\,
            in3 => \N__23115\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            clk => \N__52465\,
            ce => 'H',
            sr => \N__51995\
        );

    \current_shift_inst.PI_CTRL.error_control_30_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23112\,
            in2 => \_gnd_net_\,
            in3 => \N__23103\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_30\,
            clk => \N__52465\,
            ce => 'H',
            sr => \N__51995\
        );

    \current_shift_inst.PI_CTRL.error_control_31_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23100\,
            in2 => \_gnd_net_\,
            in3 => \N__23091\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52465\,
            ce => 'H',
            sr => \N__51995\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23087\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52459\,
            ce => 'H',
            sr => \N__52001\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23060\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52459\,
            ce => 'H',
            sr => \N__52001\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23318\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52459\,
            ce => 'H',
            sr => \N__52001\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23298\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52455\,
            ce => 'H',
            sr => \N__52009\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23279\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52455\,
            ce => 'H',
            sr => \N__52009\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23255\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52455\,
            ce => 'H',
            sr => \N__52009\
        );

    \current_shift_inst.PI_CTRL.prop_term_29_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23231\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52455\,
            ce => 'H',
            sr => \N__52009\
        );

    \current_shift_inst.PI_CTRL.prop_term_27_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23207\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52450\,
            ce => 'H',
            sr => \N__52017\
        );

    \phase_controller_inst1.start_flag_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011111000"
        )
    port map (
            in0 => \N__36588\,
            in1 => \N__36529\,
            in2 => \N__36512\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.start_flagZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52450\,
            ce => 'H',
            sr => \N__52017\
        );

    \phase_controller_inst1.state_4_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__36530\,
            in1 => \N__36589\,
            in2 => \_gnd_net_\,
            in3 => \N__36505\,
            lcout => \phase_controller_inst1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52450\,
            ce => 'H',
            sr => \N__52017\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23183\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52450\,
            ce => 'H',
            sr => \N__52017\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23516\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52442\,
            ce => 'H',
            sr => \N__52025\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23489\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52442\,
            ce => 'H',
            sr => \N__52025\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23459\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52436\,
            ce => 'H',
            sr => \N__52032\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23435\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52436\,
            ce => 'H',
            sr => \N__52032\
        );

    \current_shift_inst.PI_CTRL.prop_term_31_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23415\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52431\,
            ce => 'H',
            sr => \N__52036\
        );

    \current_shift_inst.PI_CTRL.prop_term_26_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23399\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52425\,
            ce => 'H',
            sr => \N__52041\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23378\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52425\,
            ce => 'H',
            sr => \N__52041\
        );

    \current_shift_inst.PI_CTRL.prop_term_30_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23354\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52420\,
            ce => 'H',
            sr => \N__52044\
        );

    \delay_measurement_inst.start_timer_hc_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42402\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23328\,
            ce => 'H',
            sr => \N__52046\
        );

    \delay_measurement_inst.stop_timer_hc_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42403\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23328\,
            ce => 'H',
            sr => \N__52046\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23618\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52472\,
            ce => 'H',
            sr => \N__51971\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__24276\,
            in1 => \N__24810\,
            in2 => \_gnd_net_\,
            in3 => \N__24534\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__24099\,
            in1 => \N__24840\,
            in2 => \_gnd_net_\,
            in3 => \N__24533\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__24759\,
            in1 => \N__24240\,
            in2 => \_gnd_net_\,
            in3 => \N__24535\,
            lcout => \current_shift_inst.control_input_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34236\,
            in1 => \N__32106\,
            in2 => \N__34786\,
            in3 => \N__29826\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__24536\,
            in1 => \N__25113\,
            in2 => \_gnd_net_\,
            in3 => \N__24297\,
            lcout => \current_shift_inst.control_input_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__24558\,
            in1 => \N__24357\,
            in2 => \_gnd_net_\,
            in3 => \N__24936\,
            lcout => \current_shift_inst.control_input_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001101010011"
        )
    port map (
            in0 => \N__24204\,
            in1 => \N__25011\,
            in2 => \N__24580\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__24231\,
            in1 => \N__24540\,
            in2 => \_gnd_net_\,
            in3 => \N__24732\,
            lcout => \current_shift_inst.control_input_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23778\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52443\,
            ce => 'H',
            sr => \N__51996\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23748\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52443\,
            ce => 'H',
            sr => \N__51996\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23724\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52443\,
            ce => 'H',
            sr => \N__51996\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__34787\,
            in1 => \N__34258\,
            in2 => \N__32352\,
            in3 => \N__29576\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__24475\,
            in1 => \N__24219\,
            in2 => \_gnd_net_\,
            in3 => \N__25026\,
            lcout => \current_shift_inst.control_input_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__24455\,
            in1 => \N__24705\,
            in2 => \_gnd_net_\,
            in3 => \N__24018\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__24033\,
            in1 => \N__24717\,
            in2 => \_gnd_net_\,
            in3 => \N__24454\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__24456\,
            in1 => \N__24177\,
            in2 => \_gnd_net_\,
            in3 => \N__24678\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__24666\,
            in1 => \N__24162\,
            in2 => \_gnd_net_\,
            in3 => \N__24457\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__24458\,
            in1 => \N__24396\,
            in2 => \_gnd_net_\,
            in3 => \N__24978\,
            lcout => \current_shift_inst.control_input_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37041\,
            in2 => \_gnd_net_\,
            in3 => \N__36970\,
            lcout => \phase_controller_inst1.stoper_tr.un4_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__34259\,
            in1 => \N__29921\,
            in2 => \N__34851\,
            in3 => \N__32204\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23916\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52426\,
            ce => 'H',
            sr => \N__52018\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23886\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52426\,
            ce => 'H',
            sr => \N__52018\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23862\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52426\,
            ce => 'H',
            sr => \N__52018\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23838\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52426\,
            ce => 'H',
            sr => \N__52018\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23808\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52426\,
            ce => 'H',
            sr => \N__52018\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34242\,
            in1 => \N__27293\,
            in2 => \N__34848\,
            in3 => \N__29499\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34243\,
            in1 => \N__27677\,
            in2 => \N__34847\,
            in3 => \N__29742\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34260\,
            in1 => \N__34772\,
            in2 => \N__27227\,
            in3 => \N__29457\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111000101"
        )
    port map (
            in0 => \N__27608\,
            in1 => \N__29700\,
            in2 => \N__34266\,
            in3 => \N__34773\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__34774\,
            in1 => \N__34264\,
            in2 => \N__29580\,
            in3 => \N__32345\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_28_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23991\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52409\,
            ce => 'H',
            sr => \N__52037\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__44428\,
            in1 => \N__42413\,
            in2 => \_gnd_net_\,
            in3 => \N__44335\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52409\,
            ce => 'H',
            sr => \N__52037\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52634\,
            lcout => pwm_duty_input_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52404\,
            ce => 'H',
            sr => \N__52042\
        );

    \phase_controller_inst2.state_2_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__28061\,
            in1 => \N__25841\,
            in2 => \N__23957\,
            in3 => \N__25802\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52496\,
            ce => 'H',
            sr => \N__51941\
        );

    \phase_controller_inst2.start_timer_hc_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011111000"
        )
    port map (
            in0 => \N__23950\,
            in1 => \N__25840\,
            in2 => \N__32797\,
            in3 => \N__25801\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52496\,
            ce => 'H',
            sr => \N__51941\
        );

    \phase_controller_inst2.state_1_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__25272\,
            in1 => \N__28062\,
            in2 => \N__25803\,
            in3 => \N__25240\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52496\,
            ce => 'H',
            sr => \N__51941\
        );

    \phase_controller_inst2.state_RNO_0_3_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000111111"
        )
    port map (
            in0 => \N__23961\,
            in1 => \N__25196\,
            in2 => \N__25218\,
            in3 => \N__25831\,
            lcout => \phase_controller_inst2.state_ns_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_flag_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011111000"
        )
    port map (
            in0 => \N__36565\,
            in1 => \N__24070\,
            in2 => \N__24059\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.start_flagZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52487\,
            ce => 'H',
            sr => \N__51947\
        );

    \phase_controller_inst2.state_4_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100010011000100"
        )
    port map (
            in0 => \N__36567\,
            in1 => \N__24072\,
            in2 => \N__24060\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52487\,
            ce => 'H',
            sr => \N__51947\
        );

    \phase_controller_inst2.state_3_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100011111111"
        )
    port map (
            in0 => \N__36566\,
            in1 => \N__24071\,
            in2 => \N__24058\,
            in3 => \N__24039\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52487\,
            ce => 'H',
            sr => \N__51947\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25062\,
            in2 => \N__25344\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29879\,
            in1 => \N__25656\,
            in2 => \N__25164\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34446\,
            in2 => \N__26424\,
            in3 => \N__29880\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25350\,
            in2 => \N__34637\,
            in3 => \N__24021\,
            lcout => \current_shift_inst.un38_control_input_0_s0_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34450\,
            in2 => \N__26358\,
            in3 => \N__24006\,
            lcout => \current_shift_inst.un38_control_input_0_s0_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25176\,
            in2 => \N__34638\,
            in3 => \N__24180\,
            lcout => \current_shift_inst.un38_control_input_0_s0_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34454\,
            in2 => \N__25386\,
            in3 => \N__24165\,
            lcout => \current_shift_inst.un38_control_input_0_s0_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25155\,
            in2 => \N__34639\,
            in3 => \N__24150\,
            lcout => \current_shift_inst.un38_control_input_0_s0_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34458\,
            in2 => \N__26316\,
            in3 => \N__24138\,
            lcout => \current_shift_inst.un38_control_input_0_s0_8\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25329\,
            in2 => \N__34640\,
            in3 => \N__24126\,
            lcout => \current_shift_inst.un38_control_input_0_s0_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34462\,
            in2 => \N__25323\,
            in3 => \N__24114\,
            lcout => \current_shift_inst.un38_control_input_0_s0_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25314\,
            in2 => \N__34641\,
            in3 => \N__24102\,
            lcout => \current_shift_inst.un38_control_input_0_s0_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34466\,
            in2 => \N__25308\,
            in3 => \N__24093\,
            lcout => \current_shift_inst.un38_control_input_0_s0_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25170\,
            in2 => \N__34642\,
            in3 => \N__24075\,
            lcout => \current_shift_inst.un38_control_input_0_s0_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34470\,
            in2 => \N__26340\,
            in3 => \N__24270\,
            lcout => \current_shift_inst.un38_control_input_0_s0_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28569\,
            in2 => \N__34643\,
            in3 => \N__24255\,
            lcout => \current_shift_inst.un38_control_input_0_s0_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34580\,
            in2 => \N__25443\,
            in3 => \N__24243\,
            lcout => \current_shift_inst.un38_control_input_0_s0_16\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25335\,
            in2 => \N__34743\,
            in3 => \N__24234\,
            lcout => \current_shift_inst.un38_control_input_0_s0_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34584\,
            in2 => \N__25299\,
            in3 => \N__24222\,
            lcout => \current_shift_inst.un38_control_input_0_s0_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25431\,
            in2 => \N__34744\,
            in3 => \N__24207\,
            lcout => \current_shift_inst.un38_control_input_0_s0_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34588\,
            in2 => \N__26520\,
            in3 => \N__24195\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25290\,
            in2 => \N__34745\,
            in3 => \N__24183\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34592\,
            in2 => \N__24405\,
            in3 => \N__24384\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25563\,
            in2 => \N__34746\,
            in3 => \N__24372\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34613\,
            in2 => \N__24369\,
            in3 => \N__24351\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25404\,
            in2 => \N__34763\,
            in3 => \N__24339\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34617\,
            in2 => \N__26583\,
            in3 => \N__24327\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26325\,
            in2 => \N__34764\,
            in3 => \N__24312\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34621\,
            in2 => \N__25425\,
            in3 => \N__24300\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25503\,
            in2 => \N__34765\,
            in3 => \N__24291\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25509\,
            in2 => \N__34785\,
            in3 => \N__24420\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__29031\,
            in1 => \N__25077\,
            in2 => \N__24579\,
            in3 => \N__24417\,
            lcout => \current_shift_inst.control_input_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29012\,
            in2 => \N__29881\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46342\,
            in2 => \N__25371\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46346\,
            in2 => \N__26436\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46343\,
            in2 => \N__26478\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46347\,
            in2 => \N__26448\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46344\,
            in2 => \N__26463\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46348\,
            in2 => \N__25413\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46345\,
            in2 => \N__25359\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46361\,
            in2 => \N__26532\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25497\,
            in2 => \N__46481\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46349\,
            in2 => \N__26490\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25449\,
            in2 => \N__46478\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46353\,
            in2 => \N__25458\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25491\,
            in2 => \N__46479\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46357\,
            in2 => \N__26502\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25464\,
            in2 => \N__46480\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25485\,
            in2 => \N__46482\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46368\,
            in2 => \N__25536\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25551\,
            in2 => \N__46483\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46372\,
            in2 => \N__25545\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25575\,
            in2 => \N__46484\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46376\,
            in2 => \N__25527\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25569\,
            in2 => \N__46485\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46380\,
            in2 => \N__25584\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46381\,
            in2 => \N__26673\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25608\,
            in2 => \N__46486\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46385\,
            in2 => \N__26568\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26661\,
            in2 => \N__46487\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46389\,
            in2 => \N__25680\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25686\,
            in2 => \N__46488\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46393\,
            in2 => \N__33711\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34254\,
            in2 => \_gnd_net_\,
            in3 => \N__24597\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25058\,
            in2 => \N__26399\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25661\,
            in2 => \N__25632\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34538\,
            in2 => \N__25617\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25398\,
            in2 => \N__34733\,
            in3 => \N__24708\,
            lcout => \current_shift_inst.un38_control_input_0_s1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34542\,
            in2 => \N__26610\,
            in3 => \N__24696\,
            lcout => \current_shift_inst.un38_control_input_0_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25623\,
            in2 => \N__34734\,
            in3 => \N__24681\,
            lcout => \current_shift_inst.un38_control_input_0_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34546\,
            in2 => \N__25518\,
            in3 => \N__24669\,
            lcout => \current_shift_inst.un38_control_input_0_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26373\,
            in2 => \N__34735\,
            in3 => \N__24657\,
            lcout => \current_shift_inst.un38_control_input_0_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34550\,
            in2 => \N__33393\,
            in3 => \N__24642\,
            lcout => \current_shift_inst.un38_control_input_0_s1_8\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34551\,
            in2 => \N__25602\,
            in3 => \N__24624\,
            lcout => \current_shift_inst.un38_control_input_0_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24621\,
            in2 => \N__34736\,
            in3 => \N__24600\,
            lcout => \current_shift_inst.un38_control_input_0_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34555\,
            in2 => \N__24867\,
            in3 => \N__24843\,
            lcout => \current_shift_inst.un38_control_input_0_s1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33612\,
            in2 => \N__34737\,
            in3 => \N__24828\,
            lcout => \current_shift_inst.un38_control_input_0_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34559\,
            in2 => \N__33207\,
            in3 => \N__24813\,
            lcout => \current_shift_inst.un38_control_input_0_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26544\,
            in2 => \N__34738\,
            in3 => \N__24795\,
            lcout => \current_shift_inst.un38_control_input_0_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34563\,
            in2 => \N__33303\,
            in3 => \N__24777\,
            lcout => \current_shift_inst.un38_control_input_0_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34564\,
            in2 => \N__25479\,
            in3 => \N__24762\,
            lcout => \current_shift_inst.un38_control_input_0_s1_16\,
            ltout => OPEN,
            carryin => \bfn_8_21_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26556\,
            in2 => \N__34739\,
            in3 => \N__24744\,
            lcout => \current_shift_inst.un38_control_input_0_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34568\,
            in2 => \N__24741\,
            in3 => \N__24720\,
            lcout => \current_shift_inst.un38_control_input_0_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25035\,
            in2 => \N__34740\,
            in3 => \N__25014\,
            lcout => \current_shift_inst.un38_control_input_0_s1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34572\,
            in2 => \N__26625\,
            in3 => \N__24999\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27027\,
            in2 => \N__34741\,
            in3 => \N__24981\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34576\,
            in2 => \N__29799\,
            in3 => \N__24966\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33861\,
            in2 => \N__34742\,
            in3 => \N__24945\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24942\,
            in2 => \N__34843\,
            in3 => \N__24924\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_8_22_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34750\,
            in2 => \N__26598\,
            in3 => \N__24906\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33492\,
            in2 => \N__34844\,
            in3 => \N__24885\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34754\,
            in2 => \N__26640\,
            in3 => \N__25149\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26652\,
            in2 => \N__34845\,
            in3 => \N__25131\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34758\,
            in2 => \N__25128\,
            in3 => \N__25101\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29838\,
            in2 => \N__34846\,
            in3 => \N__25083\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__34265\,
            in1 => \N__34762\,
            in2 => \_gnd_net_\,
            in3 => \N__25080\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__46489\,
            in1 => \N__25980\,
            in2 => \_gnd_net_\,
            in3 => \N__29019\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__26400\,
            in1 => \_gnd_net_\,
            in2 => \N__25065\,
            in3 => \N__46490\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S2_LC_8_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25284\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52387\,
            ce => 'H',
            sr => \N__52047\
        );

    \phase_controller_inst2.start_timer_tr_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101111111001100"
        )
    port map (
            in0 => \N__25241\,
            in1 => \N__25779\,
            in2 => \N__25280\,
            in3 => \N__28033\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52493\,
            ce => 'H',
            sr => \N__51935\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28028\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52488\,
            ce => 'H',
            sr => \N__51942\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011100000"
        )
    port map (
            in0 => \N__25216\,
            in1 => \N__27990\,
            in2 => \N__25185\,
            in3 => \N__28731\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52488\,
            ce => 'H',
            sr => \N__51942\
        );

    \phase_controller_inst2.state_0_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__25273\,
            in1 => \N__25248\,
            in2 => \N__25200\,
            in3 => \N__25217\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52488\,
            ce => 'H',
            sr => \N__51942\
        );

    \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28766\,
            in2 => \_gnd_net_\,
            in3 => \N__28034\,
            lcout => \phase_controller_inst2.stoper_tr.un4_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28776\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__28416\,
            in1 => \N__28396\,
            in2 => \_gnd_net_\,
            in3 => \N__28378\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34065\,
            in1 => \N__34491\,
            in2 => \N__26865\,
            in3 => \N__29159\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34067\,
            in1 => \N__34493\,
            in2 => \N__33255\,
            in3 => \N__33285\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__33161\,
            in1 => \N__34063\,
            in2 => \N__29310\,
            in3 => \N__25657\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34066\,
            in1 => \N__34492\,
            in2 => \N__26739\,
            in3 => \N__29088\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__34490\,
            in1 => \N__34064\,
            in2 => \N__29238\,
            in3 => \N__26976\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__34062\,
            in1 => \N__26409\,
            in2 => \_gnd_net_\,
            in3 => \N__28809\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34077\,
            in1 => \N__27738\,
            in2 => \N__34793\,
            in3 => \N__29778\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34073\,
            in1 => \N__27354\,
            in2 => \N__34791\,
            in3 => \N__29535\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__29498\,
            in1 => \N__34676\,
            in2 => \N__27294\,
            in3 => \N__34074\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34075\,
            in1 => \N__34681\,
            in2 => \N__27228\,
            in3 => \N__29456\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__33642\,
            in1 => \N__34677\,
            in2 => \N__33690\,
            in3 => \N__34076\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34078\,
            in1 => \N__27678\,
            in2 => \N__34792\,
            in3 => \N__29738\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__34683\,
            in1 => \N__34088\,
            in2 => \N__27489\,
            in3 => \N__29618\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34086\,
            in1 => \N__34685\,
            in2 => \N__32157\,
            in3 => \N__29361\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34087\,
            in1 => \N__34684\,
            in2 => \N__27612\,
            in3 => \N__29699\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__34682\,
            in1 => \N__34089\,
            in2 => \N__33600\,
            in3 => \N__29952\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28944\,
            in1 => \N__26799\,
            in2 => \_gnd_net_\,
            in3 => \N__29113\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__32301\,
            in1 => \N__34135\,
            in2 => \N__30030\,
            in3 => \N__34799\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34133\,
            in1 => \N__26972\,
            in2 => \N__34852\,
            in3 => \N__29231\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__29114\,
            in1 => \N__34134\,
            in2 => \N__26805\,
            in3 => \N__34797\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__28943\,
            in1 => \N__29299\,
            in2 => \_gnd_net_\,
            in3 => \N__33154\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__26730\,
            in1 => \N__28945\,
            in2 => \_gnd_net_\,
            in3 => \N__29083\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \N__34800\,
            in1 => \N__34235\,
            in2 => \N__29889\,
            in3 => \N__33729\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34234\,
            in1 => \N__34798\,
            in2 => \N__32211\,
            in3 => \N__29922\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28946\,
            in1 => \N__27346\,
            in2 => \_gnd_net_\,
            in3 => \N__29527\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__33241\,
            in1 => \N__33280\,
            in2 => \_gnd_net_\,
            in3 => \N__28949\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__28951\,
            in1 => \N__29356\,
            in2 => \_gnd_net_\,
            in3 => \N__32149\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__34229\,
            in1 => \N__29357\,
            in2 => \N__34853\,
            in3 => \N__32150\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__33328\,
            in1 => \N__28950\,
            in2 => \_gnd_net_\,
            in3 => \N__33367\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28948\,
            in1 => \N__33682\,
            in2 => \_gnd_net_\,
            in3 => \N__33637\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__27226\,
            in1 => \N__28947\,
            in2 => \_gnd_net_\,
            in3 => \N__29446\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__33916\,
            in1 => \N__28958\,
            in2 => \_gnd_net_\,
            in3 => \N__33880\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28956\,
            in1 => \N__27546\,
            in2 => \_gnd_net_\,
            in3 => \N__29650\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__29822\,
            in1 => \N__28957\,
            in2 => \_gnd_net_\,
            in3 => \N__32102\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__33881\,
            in1 => \N__34230\,
            in2 => \N__34854\,
            in3 => \N__33917\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28953\,
            in1 => \N__27673\,
            in2 => \_gnd_net_\,
            in3 => \N__29731\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28955\,
            in1 => \N__27604\,
            in2 => \_gnd_net_\,
            in3 => \N__29689\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28952\,
            in1 => \N__27734\,
            in2 => \_gnd_net_\,
            in3 => \N__29774\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__27482\,
            in1 => \N__29611\,
            in2 => \_gnd_net_\,
            in3 => \N__28954\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__34809\,
            in1 => \N__34195\,
            in2 => \N__26803\,
            in3 => \N__29118\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__34191\,
            in1 => \N__29917\,
            in2 => \_gnd_net_\,
            in3 => \N__32197\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__33589\,
            in1 => \N__34190\,
            in2 => \_gnd_net_\,
            in3 => \N__29945\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__34192\,
            in1 => \N__29309\,
            in2 => \N__25671\,
            in3 => \N__33162\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__34808\,
            in1 => \N__34194\,
            in2 => \N__29160\,
            in3 => \N__26861\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34193\,
            in1 => \N__34810\,
            in2 => \N__27015\,
            in3 => \N__29274\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32293\,
            in1 => \N__34189\,
            in2 => \_gnd_net_\,
            in3 => \N__30023\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34196\,
            in1 => \N__34807\,
            in2 => \N__27353\,
            in3 => \N__29534\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25969\,
            in1 => \N__28828\,
            in2 => \_gnd_net_\,
            in3 => \N__25590\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__52415\,
            ce => \N__32610\,
            sr => \N__52002\
        );

    \current_shift_inst.timer_s1.counter_1_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25957\,
            in1 => \N__33181\,
            in2 => \_gnd_net_\,
            in3 => \N__25587\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__52415\,
            ce => \N__32610\,
            sr => \N__52002\
        );

    \current_shift_inst.timer_s1.counter_2_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25970\,
            in1 => \N__26939\,
            in2 => \_gnd_net_\,
            in3 => \N__25713\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__52415\,
            ce => \N__32610\,
            sr => \N__52002\
        );

    \current_shift_inst.timer_s1.counter_3_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25958\,
            in1 => \N__26885\,
            in2 => \_gnd_net_\,
            in3 => \N__25710\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__52415\,
            ce => \N__32610\,
            sr => \N__52002\
        );

    \current_shift_inst.timer_s1.counter_4_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25971\,
            in1 => \N__26825\,
            in2 => \_gnd_net_\,
            in3 => \N__25707\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__52415\,
            ce => \N__32610\,
            sr => \N__52002\
        );

    \current_shift_inst.timer_s1.counter_5_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25959\,
            in1 => \N__26759\,
            in2 => \_gnd_net_\,
            in3 => \N__25704\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__52415\,
            ce => \N__32610\,
            sr => \N__52002\
        );

    \current_shift_inst.timer_s1.counter_6_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25972\,
            in1 => \N__26696\,
            in2 => \_gnd_net_\,
            in3 => \N__25701\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__52415\,
            ce => \N__32610\,
            sr => \N__52002\
        );

    \current_shift_inst.timer_s1.counter_7_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25960\,
            in1 => \N__27374\,
            in2 => \_gnd_net_\,
            in3 => \N__25698\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__52415\,
            ce => \N__32610\,
            sr => \N__52002\
        );

    \current_shift_inst.timer_s1.counter_8_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25956\,
            in1 => \N__27314\,
            in2 => \_gnd_net_\,
            in3 => \N__25695\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__52410\,
            ce => \N__32609\,
            sr => \N__52010\
        );

    \current_shift_inst.timer_s1.counter_9_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25968\,
            in1 => \N__27248\,
            in2 => \_gnd_net_\,
            in3 => \N__25692\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__52410\,
            ce => \N__32609\,
            sr => \N__52010\
        );

    \current_shift_inst.timer_s1.counter_10_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25953\,
            in1 => \N__27179\,
            in2 => \_gnd_net_\,
            in3 => \N__25689\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__52410\,
            ce => \N__32609\,
            sr => \N__52010\
        );

    \current_shift_inst.timer_s1.counter_11_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25965\,
            in1 => \N__27155\,
            in2 => \_gnd_net_\,
            in3 => \N__25740\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__52410\,
            ce => \N__32609\,
            sr => \N__52010\
        );

    \current_shift_inst.timer_s1.counter_12_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25954\,
            in1 => \N__27131\,
            in2 => \_gnd_net_\,
            in3 => \N__25737\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__52410\,
            ce => \N__32609\,
            sr => \N__52010\
        );

    \current_shift_inst.timer_s1.counter_13_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25966\,
            in1 => \N__27074\,
            in2 => \_gnd_net_\,
            in3 => \N__25734\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__52410\,
            ce => \N__32609\,
            sr => \N__52010\
        );

    \current_shift_inst.timer_s1.counter_14_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25955\,
            in1 => \N__27050\,
            in2 => \_gnd_net_\,
            in3 => \N__25731\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__52410\,
            ce => \N__32609\,
            sr => \N__52010\
        );

    \current_shift_inst.timer_s1.counter_15_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25967\,
            in1 => \N__27758\,
            in2 => \_gnd_net_\,
            in3 => \N__25728\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__52410\,
            ce => \N__32609\,
            sr => \N__52010\
        );

    \current_shift_inst.timer_s1.counter_16_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25944\,
            in1 => \N__27698\,
            in2 => \_gnd_net_\,
            in3 => \N__25725\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__52405\,
            ce => \N__32598\,
            sr => \N__52019\
        );

    \current_shift_inst.timer_s1.counter_17_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25961\,
            in1 => \N__27632\,
            in2 => \_gnd_net_\,
            in3 => \N__25722\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__52405\,
            ce => \N__32598\,
            sr => \N__52019\
        );

    \current_shift_inst.timer_s1.counter_18_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25945\,
            in1 => \N__27566\,
            in2 => \_gnd_net_\,
            in3 => \N__25719\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__52405\,
            ce => \N__32598\,
            sr => \N__52019\
        );

    \current_shift_inst.timer_s1.counter_19_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25962\,
            in1 => \N__27509\,
            in2 => \_gnd_net_\,
            in3 => \N__25716\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__52405\,
            ce => \N__32598\,
            sr => \N__52019\
        );

    \current_shift_inst.timer_s1.counter_20_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25946\,
            in1 => \N__27446\,
            in2 => \_gnd_net_\,
            in3 => \N__25770\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__52405\,
            ce => \N__32598\,
            sr => \N__52019\
        );

    \current_shift_inst.timer_s1.counter_21_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25963\,
            in1 => \N__27422\,
            in2 => \_gnd_net_\,
            in3 => \N__25767\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__52405\,
            ce => \N__32598\,
            sr => \N__52019\
        );

    \current_shift_inst.timer_s1.counter_22_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25947\,
            in1 => \N__27398\,
            in2 => \_gnd_net_\,
            in3 => \N__25764\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__52405\,
            ce => \N__32598\,
            sr => \N__52019\
        );

    \current_shift_inst.timer_s1.counter_23_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25964\,
            in1 => \N__27905\,
            in2 => \_gnd_net_\,
            in3 => \N__25761\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__52405\,
            ce => \N__32598\,
            sr => \N__52019\
        );

    \current_shift_inst.timer_s1.counter_24_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25931\,
            in1 => \N__27881\,
            in2 => \_gnd_net_\,
            in3 => \N__25758\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__52400\,
            ce => \N__32602\,
            sr => \N__52026\
        );

    \current_shift_inst.timer_s1.counter_25_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25973\,
            in1 => \N__27857\,
            in2 => \_gnd_net_\,
            in3 => \N__25755\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__52400\,
            ce => \N__32602\,
            sr => \N__52026\
        );

    \current_shift_inst.timer_s1.counter_26_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25932\,
            in1 => \N__27821\,
            in2 => \_gnd_net_\,
            in3 => \N__25752\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__52400\,
            ce => \N__32602\,
            sr => \N__52026\
        );

    \current_shift_inst.timer_s1.counter_27_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25974\,
            in1 => \N__27785\,
            in2 => \_gnd_net_\,
            in3 => \N__25749\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__52400\,
            ce => \N__32602\,
            sr => \N__52026\
        );

    \current_shift_inst.timer_s1.counter_28_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25933\,
            in1 => \N__27834\,
            in2 => \_gnd_net_\,
            in3 => \N__25746\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__52400\,
            ce => \N__32602\,
            sr => \N__52026\
        );

    \current_shift_inst.timer_s1.counter_29_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__27798\,
            in1 => \N__25934\,
            in2 => \_gnd_net_\,
            in3 => \N__25743\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52400\,
            ce => \N__32602\,
            sr => \N__52026\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28981\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52396\,
            ce => \N__33754\,
            sr => \N__52033\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33529\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40929\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S1_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25845\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52379\,
            ce => 'H',
            sr => \N__52048\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25797\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28051\,
            lcout => \phase_controller_inst2.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__28027\,
            in1 => \N__52083\,
            in2 => \_gnd_net_\,
            in3 => \N__28765\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32802\,
            in2 => \_gnd_net_\,
            in3 => \N__38215\,
            lcout => \phase_controller_inst2.stoper_hc.un4_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.counter_0_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26284\,
            in1 => \N__27969\,
            in2 => \N__28703\,
            in3 => \N__28704\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_7_0_\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_0\,
            clk => \N__52473\,
            ce => \N__26166\,
            sr => \N__51939\
        );

    \phase_controller_inst2.stoper_tr.counter_1_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26292\,
            in1 => \N__27948\,
            in2 => \_gnd_net_\,
            in3 => \N__25773\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_1\,
            clk => \N__52473\,
            ce => \N__26166\,
            sr => \N__51939\
        );

    \phase_controller_inst2.stoper_tr.counter_2_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26285\,
            in1 => \N__27927\,
            in2 => \_gnd_net_\,
            in3 => \N__26007\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_2\,
            clk => \N__52473\,
            ce => \N__26166\,
            sr => \N__51939\
        );

    \phase_controller_inst2.stoper_tr.counter_3_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26293\,
            in1 => \N__28251\,
            in2 => \_gnd_net_\,
            in3 => \N__26004\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_3\,
            clk => \N__52473\,
            ce => \N__26166\,
            sr => \N__51939\
        );

    \phase_controller_inst2.stoper_tr.counter_4_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26286\,
            in1 => \N__28230\,
            in2 => \_gnd_net_\,
            in3 => \N__26001\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_4\,
            clk => \N__52473\,
            ce => \N__26166\,
            sr => \N__51939\
        );

    \phase_controller_inst2.stoper_tr.counter_5_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26294\,
            in1 => \N__28209\,
            in2 => \_gnd_net_\,
            in3 => \N__25998\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_5\,
            clk => \N__52473\,
            ce => \N__26166\,
            sr => \N__51939\
        );

    \phase_controller_inst2.stoper_tr.counter_6_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26287\,
            in1 => \N__28188\,
            in2 => \_gnd_net_\,
            in3 => \N__25995\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_6\,
            clk => \N__52473\,
            ce => \N__26166\,
            sr => \N__51939\
        );

    \phase_controller_inst2.stoper_tr.counter_7_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26295\,
            in1 => \N__28167\,
            in2 => \_gnd_net_\,
            in3 => \N__25992\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_7\,
            clk => \N__52473\,
            ce => \N__26166\,
            sr => \N__51939\
        );

    \phase_controller_inst2.stoper_tr.counter_8_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26283\,
            in1 => \N__28146\,
            in2 => \_gnd_net_\,
            in3 => \N__25989\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_10_8_0_\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_8\,
            clk => \N__52466\,
            ce => \N__26167\,
            sr => \N__51943\
        );

    \phase_controller_inst2.stoper_tr.counter_9_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26291\,
            in1 => \N__28125\,
            in2 => \_gnd_net_\,
            in3 => \N__25986\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_9\,
            clk => \N__52466\,
            ce => \N__26167\,
            sr => \N__51943\
        );

    \phase_controller_inst2.stoper_tr.counter_10_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26280\,
            in1 => \N__28104\,
            in2 => \_gnd_net_\,
            in3 => \N__25983\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_10\,
            clk => \N__52466\,
            ce => \N__26167\,
            sr => \N__51943\
        );

    \phase_controller_inst2.stoper_tr.counter_11_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26288\,
            in1 => \N__28356\,
            in2 => \_gnd_net_\,
            in3 => \N__26034\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_11\,
            clk => \N__52466\,
            ce => \N__26167\,
            sr => \N__51943\
        );

    \phase_controller_inst2.stoper_tr.counter_12_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26281\,
            in1 => \N__28335\,
            in2 => \_gnd_net_\,
            in3 => \N__26031\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_12\,
            clk => \N__52466\,
            ce => \N__26167\,
            sr => \N__51943\
        );

    \phase_controller_inst2.stoper_tr.counter_13_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26289\,
            in1 => \N__28314\,
            in2 => \_gnd_net_\,
            in3 => \N__26028\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_13\,
            clk => \N__52466\,
            ce => \N__26167\,
            sr => \N__51943\
        );

    \phase_controller_inst2.stoper_tr.counter_14_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26282\,
            in1 => \N__28293\,
            in2 => \_gnd_net_\,
            in3 => \N__26025\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_14\,
            clk => \N__52466\,
            ce => \N__26167\,
            sr => \N__51943\
        );

    \phase_controller_inst2.stoper_tr.counter_15_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26290\,
            in1 => \N__28272\,
            in2 => \_gnd_net_\,
            in3 => \N__26022\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_15\,
            clk => \N__52466\,
            ce => \N__26167\,
            sr => \N__51943\
        );

    \phase_controller_inst2.stoper_tr.counter_16_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26272\,
            in1 => \N__28630\,
            in2 => \_gnd_net_\,
            in3 => \N__26019\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_16\,
            clk => \N__52461\,
            ce => \N__26168\,
            sr => \N__51945\
        );

    \phase_controller_inst2.stoper_tr.counter_17_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26276\,
            in1 => \N__28606\,
            in2 => \_gnd_net_\,
            in3 => \N__26016\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_17\,
            clk => \N__52461\,
            ce => \N__26168\,
            sr => \N__51945\
        );

    \phase_controller_inst2.stoper_tr.counter_18_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26273\,
            in1 => \N__28558\,
            in2 => \_gnd_net_\,
            in3 => \N__26013\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_18\,
            clk => \N__52461\,
            ce => \N__26168\,
            sr => \N__51945\
        );

    \phase_controller_inst2.stoper_tr.counter_19_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26277\,
            in1 => \N__28540\,
            in2 => \_gnd_net_\,
            in3 => \N__26010\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_19\,
            clk => \N__52461\,
            ce => \N__26168\,
            sr => \N__51945\
        );

    \phase_controller_inst2.stoper_tr.counter_20_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26274\,
            in1 => \N__32695\,
            in2 => \_gnd_net_\,
            in3 => \N__26061\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_20\,
            clk => \N__52461\,
            ce => \N__26168\,
            sr => \N__51945\
        );

    \phase_controller_inst2.stoper_tr.counter_21_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26278\,
            in1 => \N__32713\,
            in2 => \_gnd_net_\,
            in3 => \N__26058\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_21\,
            clk => \N__52461\,
            ce => \N__26168\,
            sr => \N__51945\
        );

    \phase_controller_inst2.stoper_tr.counter_22_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26275\,
            in1 => \N__32955\,
            in2 => \_gnd_net_\,
            in3 => \N__26055\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_22\,
            clk => \N__52461\,
            ce => \N__26168\,
            sr => \N__51945\
        );

    \phase_controller_inst2.stoper_tr.counter_23_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26279\,
            in1 => \N__32973\,
            in2 => \_gnd_net_\,
            in3 => \N__26052\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_23\,
            clk => \N__52461\,
            ce => \N__26168\,
            sr => \N__51945\
        );

    \phase_controller_inst2.stoper_tr.counter_24_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26264\,
            in1 => \N__28665\,
            in2 => \_gnd_net_\,
            in3 => \N__26049\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_24\,
            clk => \N__52457\,
            ce => \N__26169\,
            sr => \N__51951\
        );

    \phase_controller_inst2.stoper_tr.counter_25_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26268\,
            in1 => \N__28680\,
            in2 => \_gnd_net_\,
            in3 => \N__26046\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_25\,
            clk => \N__52457\,
            ce => \N__26169\,
            sr => \N__51951\
        );

    \phase_controller_inst2.stoper_tr.counter_26_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26265\,
            in1 => \N__32842\,
            in2 => \_gnd_net_\,
            in3 => \N__26043\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_26\,
            clk => \N__52457\,
            ce => \N__26169\,
            sr => \N__51951\
        );

    \phase_controller_inst2.stoper_tr.counter_27_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26269\,
            in1 => \N__32872\,
            in2 => \_gnd_net_\,
            in3 => \N__26040\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_27\,
            clk => \N__52457\,
            ce => \N__26169\,
            sr => \N__51951\
        );

    \phase_controller_inst2.stoper_tr.counter_28_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26266\,
            in1 => \N__28380\,
            in2 => \_gnd_net_\,
            in3 => \N__26037\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_28\,
            clk => \N__52457\,
            ce => \N__26169\,
            sr => \N__51951\
        );

    \phase_controller_inst2.stoper_tr.counter_29_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26270\,
            in1 => \N__28398\,
            in2 => \_gnd_net_\,
            in3 => \N__26301\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_29\,
            clk => \N__52457\,
            ce => \N__26169\,
            sr => \N__51951\
        );

    \phase_controller_inst2.stoper_tr.counter_30_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26267\,
            in1 => \N__28452\,
            in2 => \_gnd_net_\,
            in3 => \N__26298\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_29\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_30\,
            clk => \N__52457\,
            ce => \N__26169\,
            sr => \N__51951\
        );

    \phase_controller_inst2.stoper_tr.counter_31_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26271\,
            in1 => \N__28470\,
            in2 => \_gnd_net_\,
            in3 => \N__26172\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52457\,
            ce => \N__26169\,
            sr => \N__51951\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_28_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40470\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52451\,
            ce => \N__36325\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__28468\,
            in1 => \N__28450\,
            in2 => \_gnd_net_\,
            in3 => \N__28419\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26151\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52444\,
            ce => 'H',
            sr => \N__51956\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26121\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52444\,
            ce => 'H',
            sr => \N__51956\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26102\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52444\,
            ce => 'H',
            sr => \N__51956\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26081\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52444\,
            ce => 'H',
            sr => \N__51956\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28988\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52438\,
            ce => \N__33759\,
            sr => \N__51960\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__27007\,
            in1 => \N__34061\,
            in2 => \N__34860\,
            in3 => \N__29270\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29330\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34060\,
            in2 => \N__26403\,
            in3 => \N__28802\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__26735\,
            in1 => \N__34068\,
            in2 => \N__29087\,
            in3 => \N__34782\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34069\,
            in1 => \N__26918\,
            in2 => \N__34850\,
            in3 => \N__29189\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__29394\,
            in1 => \N__34784\,
            in2 => \N__27111\,
            in3 => \N__34071\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34072\,
            in1 => \N__32256\,
            in2 => \N__34849\,
            in3 => \N__29982\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__33411\,
            in1 => \N__34783\,
            in2 => \N__33452\,
            in3 => \N__34070\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26856\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26734\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28881\,
            in1 => \N__26965\,
            in2 => \_gnd_net_\,
            in3 => \N__29224\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28883\,
            in1 => \N__26857\,
            in2 => \_gnd_net_\,
            in3 => \N__29143\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26964\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28882\,
            in1 => \N__26917\,
            in2 => \_gnd_net_\,
            in3 => \N__29185\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26804\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27279\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28880\,
            in1 => \N__27014\,
            in2 => \_gnd_net_\,
            in3 => \N__29263\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33438\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34136\,
            in1 => \N__34893\,
            in2 => \N__27110\,
            in3 => \N__29390\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28908\,
            in1 => \N__33439\,
            in2 => \_gnd_net_\,
            in3 => \N__33409\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26916\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__29658\,
            in1 => \N__34137\,
            in2 => \N__34908\,
            in3 => \N__27541\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__27103\,
            in1 => \N__28910\,
            in2 => \_gnd_net_\,
            in3 => \N__29389\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__28909\,
            in1 => \_gnd_net_\,
            in2 => \N__27289\,
            in3 => \N__29482\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27006\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33231\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_0_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47157\,
            in2 => \_gnd_net_\,
            in3 => \N__47642\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52416\,
            ce => \N__43466\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27603\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27213\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27540\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33669\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27474\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__34188\,
            in1 => \N__34898\,
            in2 => \N__33513\,
            in3 => \N__33545\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27723\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34185\,
            in1 => \N__33544\,
            in2 => \_gnd_net_\,
            in3 => \N__33508\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33357\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34187\,
            in1 => \N__34897\,
            in2 => \N__27733\,
            in3 => \N__29770\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27672\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__28962\,
            in1 => \N__32338\,
            in2 => \_gnd_net_\,
            in3 => \N__29566\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32251\,
            in1 => \N__34186\,
            in2 => \_gnd_net_\,
            in3 => \N__29971\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__34901\,
            in1 => \N__34202\,
            in2 => \N__33596\,
            in3 => \N__29944\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27094\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__34899\,
            in1 => \N__34201\,
            in2 => \N__29978\,
            in3 => \N__32252\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27329\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__34903\,
            in1 => \N__34198\,
            in2 => \N__29657\,
            in3 => \N__27545\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__34197\,
            in1 => \N__34900\,
            in2 => \N__29199\,
            in3 => \N__26919\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__34904\,
            in1 => \N__34200\,
            in2 => \N__32300\,
            in3 => \N__30022\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__34199\,
            in1 => \N__34902\,
            in2 => \N__29619\,
            in3 => \N__27481\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26935\,
            in2 => \N__28832\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_10_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__52401\,
            ce => \N__33756\,
            sr => \N__51997\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26881\,
            in2 => \N__33185\,
            in3 => \N__26943\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__52401\,
            ce => \N__33756\,
            sr => \N__51997\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26821\,
            in2 => \N__26940\,
            in3 => \N__26889\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__52401\,
            ce => \N__33756\,
            sr => \N__51997\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26755\,
            in2 => \N__26886\,
            in3 => \N__26829\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__52401\,
            ce => \N__33756\,
            sr => \N__51997\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26692\,
            in2 => \N__26826\,
            in3 => \N__26763\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__52401\,
            ce => \N__33756\,
            sr => \N__51997\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27370\,
            in2 => \N__26760\,
            in3 => \N__26700\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__52401\,
            ce => \N__33756\,
            sr => \N__51997\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27310\,
            in2 => \N__26697\,
            in3 => \N__26676\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__52401\,
            ce => \N__33756\,
            sr => \N__51997\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27244\,
            in2 => \N__27375\,
            in3 => \N__27318\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__52401\,
            ce => \N__33756\,
            sr => \N__51997\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27175\,
            in2 => \N__27315\,
            in3 => \N__27252\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__52397\,
            ce => \N__33755\,
            sr => \N__52003\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27151\,
            in2 => \N__27249\,
            in3 => \N__27183\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__52397\,
            ce => \N__33755\,
            sr => \N__52003\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27127\,
            in2 => \N__27180\,
            in3 => \N__27159\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__52397\,
            ce => \N__33755\,
            sr => \N__52003\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27070\,
            in2 => \N__27156\,
            in3 => \N__27135\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__52397\,
            ce => \N__33755\,
            sr => \N__52003\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27046\,
            in2 => \N__27132\,
            in3 => \N__27078\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__52397\,
            ce => \N__33755\,
            sr => \N__52003\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27754\,
            in2 => \N__27075\,
            in3 => \N__27054\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__52397\,
            ce => \N__33755\,
            sr => \N__52003\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27694\,
            in2 => \N__27051\,
            in3 => \N__27030\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__52397\,
            ce => \N__33755\,
            sr => \N__52003\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27628\,
            in2 => \N__27759\,
            in3 => \N__27702\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__52397\,
            ce => \N__33755\,
            sr => \N__52003\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27562\,
            in2 => \N__27699\,
            in3 => \N__27636\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__52392\,
            ce => \N__33753\,
            sr => \N__52011\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27505\,
            in2 => \N__27633\,
            in3 => \N__27570\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__52392\,
            ce => \N__33753\,
            sr => \N__52011\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27442\,
            in2 => \N__27567\,
            in3 => \N__27513\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__52392\,
            ce => \N__33753\,
            sr => \N__52011\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27418\,
            in2 => \N__27510\,
            in3 => \N__27450\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__52392\,
            ce => \N__33753\,
            sr => \N__52011\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27394\,
            in2 => \N__27447\,
            in3 => \N__27426\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__52392\,
            ce => \N__33753\,
            sr => \N__52011\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27901\,
            in2 => \N__27423\,
            in3 => \N__27402\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__52392\,
            ce => \N__33753\,
            sr => \N__52011\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27877\,
            in2 => \N__27399\,
            in3 => \N__27378\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__52392\,
            ce => \N__33753\,
            sr => \N__52011\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27853\,
            in2 => \N__27906\,
            in3 => \N__27885\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__52392\,
            ce => \N__33753\,
            sr => \N__52011\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27817\,
            in2 => \N__27882\,
            in3 => \N__27861\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__52389\,
            ce => \N__33752\,
            sr => \N__52020\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27781\,
            in2 => \N__27858\,
            in3 => \N__27837\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__52389\,
            ce => \N__33752\,
            sr => \N__52020\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27833\,
            in2 => \N__27822\,
            in3 => \N__27801\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__52389\,
            ce => \N__33752\,
            sr => \N__52020\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27797\,
            in2 => \N__27786\,
            in3 => \N__27765\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__52389\,
            ce => \N__33752\,
            sr => \N__52020\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27762\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37040\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52384\,
            ce => 'H',
            sr => \N__52030\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36959\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__35787\,
            in1 => \N__34950\,
            in2 => \_gnd_net_\,
            in3 => \N__35813\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__27985\,
            in1 => \N__28029\,
            in2 => \_gnd_net_\,
            in3 => \N__28778\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__38772\,
            in1 => \N__32817\,
            in2 => \N__28071\,
            in3 => \N__28055\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52474\,
            ce => 'H',
            sr => \N__51932\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32801\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52474\,
            ce => 'H',
            sr => \N__51932\
        );

    \phase_controller_inst2.stoper_hc.running_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000101110"
        )
    port map (
            in0 => \N__32816\,
            in1 => \N__32800\,
            in2 => \N__38220\,
            in3 => \N__38771\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52474\,
            ce => 'H',
            sr => \N__51932\
        );

    \phase_controller_inst2.stoper_tr.running_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000101110"
        )
    port map (
            in0 => \N__27989\,
            in1 => \N__28035\,
            in2 => \N__28782\,
            in3 => \N__28730\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52474\,
            ce => 'H',
            sr => \N__51932\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33054\,
            in2 => \N__27957\,
            in3 => \N__27968\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32736\,
            in2 => \N__27936\,
            in3 => \N__27947\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32742\,
            in2 => \N__27915\,
            in3 => \N__27926\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28250\,
            in1 => \N__32754\,
            in2 => \N__28239\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32928\,
            in2 => \N__28218\,
            in3 => \N__28229\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32748\,
            in2 => \N__28197\,
            in3 => \N__28208\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28187\,
            in1 => \N__33009\,
            in2 => \N__28176\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36426\,
            in2 => \N__28155\,
            in3 => \N__28166\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32730\,
            in2 => \N__28134\,
            in3 => \N__28145\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32916\,
            in2 => \N__28113\,
            in3 => \N__28124\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28103\,
            in1 => \N__33066\,
            in2 => \N__28092\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33042\,
            in2 => \N__28344\,
            in3 => \N__28355\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32991\,
            in2 => \N__28323\,
            in3 => \N__28334\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28313\,
            in1 => \N__32907\,
            in2 => \N__28302\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28292\,
            in1 => \N__33480\,
            in2 => \N__28281\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36489\,
            in2 => \N__28260\,
            in3 => \N__28271\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28590\,
            in2 => \N__28644\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28581\,
            in2 => \N__28524\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32679\,
            in2 => \N__32724\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32979\,
            in2 => \N__32937\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28650\,
            in2 => \N__28428\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28509\,
            in2 => \N__33120\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28362\,
            in2 => \N__28500\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28434\,
            in2 => \N__28485\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28473\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__28418\,
            in1 => \N__28469\,
            in2 => \_gnd_net_\,
            in3 => \N__28451\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101010001"
        )
    port map (
            in0 => \N__28678\,
            in1 => \N__28663\,
            in2 => \N__33029\,
            in3 => \N__32888\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__28417\,
            in1 => \N__28397\,
            in2 => \_gnd_net_\,
            in3 => \N__28379\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28777\,
            in2 => \_gnd_net_\,
            in3 => \N__28720\,
            lcout => \phase_controller_inst2.stoper_tr.counter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__52084\,
            in1 => \N__33105\,
            in2 => \_gnd_net_\,
            in3 => \N__39209\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100010000"
        )
    port map (
            in0 => \N__28679\,
            in1 => \N__28664\,
            in2 => \N__33030\,
            in3 => \N__32889\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__36393\,
            in1 => \N__28632\,
            in2 => \N__28614\,
            in3 => \N__32898\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__36392\,
            in1 => \N__28631\,
            in2 => \N__28613\,
            in3 => \N__32897\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011011101"
        )
    port map (
            in0 => \N__28541\,
            in1 => \N__36377\,
            in2 => \N__36411\,
            in3 => \N__28559\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34079\,
            in1 => \N__33378\,
            in2 => \N__34859\,
            in3 => \N__33333\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__28560\,
            in1 => \N__36407\,
            in2 => \N__36378\,
            in3 => \N__28542\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011101111"
        )
    port map (
            in0 => \N__36477\,
            in1 => \N__36030\,
            in2 => \N__32849\,
            in3 => \N__32876\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33096\,
            in2 => \_gnd_net_\,
            in3 => \N__39197\,
            lcout => \phase_controller_inst1.stoper_hc.un4_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__29043\,
            in1 => \N__29049\,
            in2 => \N__39231\,
            in3 => \N__36783\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52433\,
            ce => 'H',
            sr => \N__51957\
        );

    \phase_controller_inst1.stoper_hc.running_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111001001110"
        )
    port map (
            in0 => \N__33095\,
            in1 => \N__29042\,
            in2 => \N__39207\,
            in3 => \N__39230\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52433\,
            ce => 'H',
            sr => \N__51957\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__29041\,
            in1 => \N__33094\,
            in2 => \_gnd_net_\,
            in3 => \N__39193\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34090\,
            in2 => \_gnd_net_\,
            in3 => \N__34775\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28800\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__28801\,
            in1 => \_gnd_net_\,
            in2 => \N__29022\,
            in3 => \N__28876\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28995\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52428\,
            ce => \N__33758\,
            sr => \N__51961\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28839\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52428\,
            ce => \N__33758\,
            sr => \N__51961\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33459\,
            in2 => \N__29334\,
            in3 => \N__29329\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29280\,
            in2 => \_gnd_net_\,
            in3 => \N__29247\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29244\,
            in2 => \_gnd_net_\,
            in3 => \N__29208\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29205\,
            in2 => \_gnd_net_\,
            in3 => \N__29169\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29166\,
            in2 => \_gnd_net_\,
            in3 => \N__29127\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29124\,
            in2 => \_gnd_net_\,
            in3 => \N__29097\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29094\,
            in2 => \_gnd_net_\,
            in3 => \N__29061\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29058\,
            in2 => \_gnd_net_\,
            in3 => \N__29052\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29547\,
            in3 => \N__29508\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29505\,
            in2 => \_gnd_net_\,
            in3 => \N__29466\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29463\,
            in2 => \_gnd_net_\,
            in3 => \N__29424\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29421\,
            in2 => \_gnd_net_\,
            in3 => \N__29415\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29412\,
            in2 => \_gnd_net_\,
            in3 => \N__29406\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29403\,
            in2 => \_gnd_net_\,
            in3 => \N__29376\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29373\,
            in2 => \_gnd_net_\,
            in3 => \N__29364\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32121\,
            in2 => \_gnd_net_\,
            in3 => \N__29337\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29784\,
            in2 => \_gnd_net_\,
            in3 => \N__29751\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29748\,
            in2 => \_gnd_net_\,
            in3 => \N__29709\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29706\,
            in2 => \_gnd_net_\,
            in3 => \N__29667\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29664\,
            in2 => \_gnd_net_\,
            in3 => \N__29628\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29625\,
            in2 => \_gnd_net_\,
            in3 => \N__29589\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32064\,
            in2 => \_gnd_net_\,
            in3 => \N__29586\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33696\,
            in2 => \_gnd_net_\,
            in3 => \N__29583\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32310\,
            in2 => \_gnd_net_\,
            in3 => \N__29550\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32265\,
            in2 => \_gnd_net_\,
            in3 => \N__30003\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30000\,
            in2 => \_gnd_net_\,
            in3 => \N__29985\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32223\,
            in2 => \_gnd_net_\,
            in3 => \N__29955\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33555\,
            in2 => \_gnd_net_\,
            in3 => \N__29925\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32166\,
            in2 => \_gnd_net_\,
            in3 => \N__29895\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29892\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \N__29888\,
            in1 => \N__34887\,
            in2 => \N__29841\,
            in3 => \N__34238\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34237\,
            in1 => \N__32098\,
            in2 => \N__34905\,
            in3 => \N__29818\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36729\,
            in2 => \N__36708\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30435\,
            in2 => \N__30408\,
            in3 => \N__30393\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__52402\,
            ce => 'H',
            sr => \N__51986\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30390\,
            in2 => \N__30375\,
            in3 => \N__30324\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__52402\,
            ce => 'H',
            sr => \N__51986\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30321\,
            in2 => \N__30309\,
            in3 => \N__30270\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__52402\,
            ce => 'H',
            sr => \N__51986\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30267\,
            in2 => \N__30252\,
            in3 => \N__30204\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__52402\,
            ce => 'H',
            sr => \N__51986\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30201\,
            in2 => \N__30186\,
            in3 => \N__30147\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__52402\,
            ce => 'H',
            sr => \N__51986\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30144\,
            in2 => \N__30129\,
            in3 => \N__30084\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__52402\,
            ce => 'H',
            sr => \N__51986\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30081\,
            in2 => \N__30072\,
            in3 => \N__30033\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__52402\,
            ce => 'H',
            sr => \N__51986\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30954\,
            in2 => \N__30942\,
            in3 => \N__30894\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__52398\,
            ce => 'H',
            sr => \N__51993\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30891\,
            in2 => \N__30873\,
            in3 => \N__30825\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__52398\,
            ce => 'H',
            sr => \N__51993\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30822\,
            in2 => \N__30807\,
            in3 => \N__30756\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__52398\,
            ce => 'H',
            sr => \N__51993\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30753\,
            in2 => \N__30738\,
            in3 => \N__30687\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__52398\,
            ce => 'H',
            sr => \N__51993\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30684\,
            in2 => \N__30669\,
            in3 => \N__30627\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__52398\,
            ce => 'H',
            sr => \N__51993\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30624\,
            in2 => \N__30609\,
            in3 => \N__30573\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__52398\,
            ce => 'H',
            sr => \N__51993\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30570\,
            in2 => \N__30555\,
            in3 => \N__30498\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__52398\,
            ce => 'H',
            sr => \N__51993\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30495\,
            in2 => \N__30483\,
            in3 => \N__30438\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__52398\,
            ce => 'H',
            sr => \N__51993\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31452\,
            in2 => \N__31443\,
            in3 => \N__31392\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_21_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__52393\,
            ce => 'H',
            sr => \N__51998\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31389\,
            in2 => \N__31374\,
            in3 => \N__31329\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__52393\,
            ce => 'H',
            sr => \N__51998\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31326\,
            in2 => \N__31308\,
            in3 => \N__31260\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__52393\,
            ce => 'H',
            sr => \N__51998\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31257\,
            in2 => \N__31242\,
            in3 => \N__31188\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__52393\,
            ce => 'H',
            sr => \N__51998\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31185\,
            in2 => \N__31173\,
            in3 => \N__31134\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__52393\,
            ce => 'H',
            sr => \N__51998\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31131\,
            in2 => \N__31119\,
            in3 => \N__31077\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__52393\,
            ce => 'H',
            sr => \N__51998\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31074\,
            in2 => \N__31062\,
            in3 => \N__31017\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__52393\,
            ce => 'H',
            sr => \N__51998\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31014\,
            in2 => \N__30999\,
            in3 => \N__30957\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__52393\,
            ce => 'H',
            sr => \N__51998\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32046\,
            in2 => \N__32028\,
            in3 => \N__31983\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__52390\,
            ce => 'H',
            sr => \N__52004\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31980\,
            in2 => \N__31965\,
            in3 => \N__31920\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__52390\,
            ce => 'H',
            sr => \N__52004\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31917\,
            in2 => \N__31899\,
            in3 => \N__31851\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__52390\,
            ce => 'H',
            sr => \N__52004\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31848\,
            in2 => \N__31839\,
            in3 => \N__31785\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__52390\,
            ce => 'H',
            sr => \N__52004\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31782\,
            in2 => \N__31764\,
            in3 => \N__31725\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__52390\,
            ce => 'H',
            sr => \N__52004\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31722\,
            in2 => \N__31713\,
            in3 => \N__31662\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__52390\,
            ce => 'H',
            sr => \N__52004\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31659\,
            in1 => \N__31488\,
            in2 => \_gnd_net_\,
            in3 => \N__31473\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52390\,
            ce => 'H',
            sr => \N__52004\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__36885\,
            in1 => \N__37036\,
            in2 => \_gnd_net_\,
            in3 => \N__36949\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32328\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32276\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32234\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32182\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32140\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__35844\,
            in1 => \N__35300\,
            in2 => \N__35876\,
            in3 => \N__35286\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32088\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32052\,
            in2 => \N__34986\,
            in3 => \N__35247\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_11_25_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35082\,
            in2 => \N__32439\,
            in3 => \N__35232\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35076\,
            in2 => \N__32430\,
            in3 => \N__35214\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35088\,
            in2 => \N__32421\,
            in3 => \N__35193\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35307\,
            in2 => \N__32412\,
            in3 => \N__35172\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35094\,
            in2 => \N__32400\,
            in3 => \N__35154\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35469\,
            in1 => \N__35070\,
            in2 => \N__32391\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33813\,
            in2 => \N__32379\,
            in3 => \N__35451\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35064\,
            in2 => \N__32370\,
            in3 => \N__35433\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_11_26_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35019\,
            in2 => \N__32361\,
            in3 => \N__35415\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33837\,
            in2 => \N__32505\,
            in3 => \N__35397\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33801\,
            in2 => \N__32496\,
            in3 => \N__35379\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33825\,
            in2 => \N__32484\,
            in3 => \N__35361\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35343\,
            in1 => \N__35058\,
            in2 => \N__32472\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35325\,
            in1 => \N__33789\,
            in2 => \N__32460\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33849\,
            in2 => \N__32448\,
            in3 => \N__35562\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37932\,
            in2 => \N__37851\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_27_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38283\,
            in2 => \N__38358\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_11_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32664\,
            in2 => \N__32652\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32658\,
            in2 => \N__32673\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32619\,
            in2 => \N__32640\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35268\,
            in2 => \N__32535\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32523\,
            in2 => \N__32514\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32628\,
            in2 => \N__32550\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32517\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36966\,
            in2 => \_gnd_net_\,
            in3 => \N__36896\,
            lcout => \phase_controller_inst1.stoper_tr.counter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__34944\,
            in1 => \N__35786\,
            in2 => \_gnd_net_\,
            in3 => \N__35814\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__33776\,
            in1 => \N__35938\,
            in2 => \N__35042\,
            in3 => \N__35485\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_11_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__35114\,
            in1 => \N__35007\,
            in2 => \N__35511\,
            in3 => \N__35531\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__33777\,
            in1 => \N__35939\,
            in2 => \N__35043\,
            in3 => \N__35486\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_11_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010111011"
        )
    port map (
            in0 => \N__35006\,
            in1 => \N__35506\,
            in2 => \N__35115\,
            in3 => \N__35530\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_11_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011110101"
        )
    port map (
            in0 => \N__35896\,
            in1 => \N__35132\,
            in2 => \N__34971\,
            in3 => \N__35920\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__35756\,
            in1 => \N__35597\,
            in2 => \_gnd_net_\,
            in3 => \N__34945\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__35133\,
            in1 => \N__34970\,
            in2 => \N__35901\,
            in3 => \N__35921\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_11_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__41171\,
            in1 => \N__40893\,
            in2 => \_gnd_net_\,
            in3 => \N__40925\,
            lcout => \current_shift_inst.timer_s1.N_154_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_11_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35755\,
            in2 => \N__34949\,
            in3 => \N__35596\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32799\,
            in2 => \N__38212\,
            in3 => \N__32815\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__52082\,
            in1 => \N__32798\,
            in2 => \_gnd_net_\,
            in3 => \N__38214\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_3_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37293\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52460\,
            ce => \N__36314\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_5_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37233\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52460\,
            ce => \N__36314\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_2_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37323\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52460\,
            ce => \N__36314\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_1_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37353\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52460\,
            ce => \N__36314\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_8_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37152\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52456\,
            ce => \N__36324\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__36462\,
            in1 => \N__32715\,
            in2 => \N__36360\,
            in3 => \N__32697\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__36461\,
            in1 => \N__32714\,
            in2 => \N__36359\,
            in3 => \N__32696\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011010100"
        )
    port map (
            in0 => \N__32972\,
            in1 => \N__36042\,
            in2 => \N__36447\,
            in3 => \N__32954\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011110101"
        )
    port map (
            in0 => \N__32971\,
            in1 => \N__36041\,
            in2 => \N__36446\,
            in3 => \N__32953\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__36098\,
            in1 => \N__36248\,
            in2 => \_gnd_net_\,
            in3 => \N__38914\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__36097\,
            in1 => \N__36247\,
            in2 => \_gnd_net_\,
            in3 => \N__38913\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_4_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37263\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52437\,
            ce => \N__36332\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_9_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37548\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52437\,
            ce => \N__36332\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_13_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37461\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52437\,
            ce => \N__36332\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_17_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37377\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52437\,
            ce => \N__36332\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_25_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37569\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52432\,
            ce => \N__36333\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__32877\,
            in1 => \N__36029\,
            in2 => \N__32850\,
            in3 => \N__36476\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33100\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52427\,
            ce => 'H',
            sr => \N__51953\
        );

    \phase_controller_inst1.state_1_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__37072\,
            in1 => \N__38246\,
            in2 => \N__36758\,
            in3 => \N__36787\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52427\,
            ce => 'H',
            sr => \N__51953\
        );

    \phase_controller_inst1.start_timer_hc_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011111000"
        )
    port map (
            in0 => \N__41217\,
            in1 => \N__36646\,
            in2 => \N__33104\,
            in3 => \N__36753\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52427\,
            ce => 'H',
            sr => \N__51953\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_10_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37524\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52421\,
            ce => \N__36334\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_0_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42297\,
            in2 => \_gnd_net_\,
            in3 => \N__39615\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52421\,
            ce => \N__36334\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_11_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37503\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52421\,
            ce => \N__36334\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_24_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37590\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52421\,
            ce => \N__36334\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_6_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37202\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52421\,
            ce => \N__36334\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_12_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37482\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52421\,
            ce => \N__36334\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_14_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37440\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52421\,
            ce => \N__36334\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36844\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33468\,
            ce => 'H',
            sr => \N__51962\
        );

    \delay_measurement_inst.start_timer_tr_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36845\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33468\,
            ce => 'H',
            sr => \N__51962\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33136\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37737\,
            in2 => \_gnd_net_\,
            in3 => \N__36817\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_157_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__34855\,
            in1 => \N__34209\,
            in2 => \N__33453\,
            in3 => \N__33410\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__34211\,
            in1 => \N__33374\,
            in2 => \N__33332\,
            in3 => \N__34857\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__34210\,
            in1 => \N__34856\,
            in2 => \N__33281\,
            in3 => \N__33248\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33189\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52406\,
            ce => \N__33757\,
            sr => \N__51972\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__34208\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33722\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33915\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34244\,
            in1 => \N__34858\,
            in2 => \N__33689\,
            in3 => \N__33638\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36759\,
            in2 => \_gnd_net_\,
            in3 => \N__36794\,
            lcout => \phase_controller_inst1.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__52085\,
            in1 => \N__37013\,
            in2 => \_gnd_net_\,
            in3 => \N__36974\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42503\,
            in2 => \_gnd_net_\,
            in3 => \N__42522\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33588\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__34907\,
            in1 => \N__34246\,
            in2 => \N__33549\,
            in3 => \N__33509\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__34906\,
            in1 => \N__34245\,
            in2 => \N__33921\,
            in3 => \N__33882\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_15_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37412\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52391\,
            ce => \N__38374\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_10_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37517\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52391\,
            ce => \N__38374\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_12_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37475\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52391\,
            ce => \N__38374\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_7_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37172\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52388\,
            ce => \N__38405\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_16_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37391\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52388\,
            ce => \N__38405\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_11_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37496\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52388\,
            ce => \N__38405\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_14_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37433\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52388\,
            ce => \N__38405\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_22_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37625\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52388\,
            ce => \N__38405\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_13_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37454\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52388\,
            ce => \N__38405\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_23_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37604\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52388\,
            ce => \N__38405\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_27_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37757\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52383\,
            ce => \N__38423\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_9_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37541\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52383\,
            ce => \N__38423\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_18_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37694\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52383\,
            ce => \N__38423\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_21_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37646\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52383\,
            ce => \N__38423\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_0_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42296\,
            in2 => \_gnd_net_\,
            in3 => \N__39614\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52380\,
            ce => \N__38409\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_25_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37562\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52380\,
            ce => \N__38409\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_28_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40463\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52380\,
            ce => \N__38409\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_17_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37373\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52380\,
            ce => \N__38409\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_26_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37778\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52380\,
            ce => \N__38409\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_24_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37583\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52380\,
            ce => \N__38409\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_20_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37676\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52376\,
            ce => \N__38404\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_5_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37229\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52376\,
            ce => \N__38404\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_3_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37289\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52376\,
            ce => \N__38404\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37352\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52373\,
            ce => \N__38419\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_2_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37319\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52373\,
            ce => \N__38419\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_6_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37203\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52373\,
            ce => \N__38419\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_8_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37148\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52373\,
            ce => \N__38419\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_4_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37262\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52373\,
            ce => \N__38419\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__35840\,
            in1 => \N__35301\,
            in2 => \N__35877\,
            in3 => \N__35285\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.counter_0_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35705\,
            in1 => \N__35246\,
            in2 => \N__35262\,
            in3 => \N__35261\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_27_0_\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_0\,
            clk => \N__52370\,
            ce => \N__35580\,
            sr => \N__52034\
        );

    \phase_controller_inst1.stoper_tr.counter_1_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35733\,
            in1 => \N__35231\,
            in2 => \_gnd_net_\,
            in3 => \N__35217\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_1\,
            clk => \N__52370\,
            ce => \N__35580\,
            sr => \N__52034\
        );

    \phase_controller_inst1.stoper_tr.counter_2_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35706\,
            in1 => \N__35210\,
            in2 => \_gnd_net_\,
            in3 => \N__35196\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_2\,
            clk => \N__52370\,
            ce => \N__35580\,
            sr => \N__52034\
        );

    \phase_controller_inst1.stoper_tr.counter_3_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35734\,
            in1 => \N__35189\,
            in2 => \_gnd_net_\,
            in3 => \N__35175\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_3\,
            clk => \N__52370\,
            ce => \N__35580\,
            sr => \N__52034\
        );

    \phase_controller_inst1.stoper_tr.counter_4_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35707\,
            in1 => \N__35171\,
            in2 => \_gnd_net_\,
            in3 => \N__35157\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_4\,
            clk => \N__52370\,
            ce => \N__35580\,
            sr => \N__52034\
        );

    \phase_controller_inst1.stoper_tr.counter_5_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35735\,
            in1 => \N__35150\,
            in2 => \_gnd_net_\,
            in3 => \N__35136\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_5\,
            clk => \N__52370\,
            ce => \N__35580\,
            sr => \N__52034\
        );

    \phase_controller_inst1.stoper_tr.counter_6_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35708\,
            in1 => \N__35468\,
            in2 => \_gnd_net_\,
            in3 => \N__35454\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_6\,
            clk => \N__52370\,
            ce => \N__35580\,
            sr => \N__52034\
        );

    \phase_controller_inst1.stoper_tr.counter_7_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35736\,
            in1 => \N__35450\,
            in2 => \_gnd_net_\,
            in3 => \N__35436\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_7\,
            clk => \N__52370\,
            ce => \N__35580\,
            sr => \N__52034\
        );

    \phase_controller_inst1.stoper_tr.counter_8_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35712\,
            in1 => \N__35432\,
            in2 => \_gnd_net_\,
            in3 => \N__35418\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_28_0_\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_8\,
            clk => \N__52367\,
            ce => \N__35579\,
            sr => \N__52038\
        );

    \phase_controller_inst1.stoper_tr.counter_9_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35729\,
            in1 => \N__35414\,
            in2 => \_gnd_net_\,
            in3 => \N__35400\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_9\,
            clk => \N__52367\,
            ce => \N__35579\,
            sr => \N__52038\
        );

    \phase_controller_inst1.stoper_tr.counter_10_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35709\,
            in1 => \N__35396\,
            in2 => \_gnd_net_\,
            in3 => \N__35382\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_10\,
            clk => \N__52367\,
            ce => \N__35579\,
            sr => \N__52038\
        );

    \phase_controller_inst1.stoper_tr.counter_11_LC_12_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35726\,
            in1 => \N__35378\,
            in2 => \_gnd_net_\,
            in3 => \N__35364\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_11\,
            clk => \N__52367\,
            ce => \N__35579\,
            sr => \N__52038\
        );

    \phase_controller_inst1.stoper_tr.counter_12_LC_12_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35710\,
            in1 => \N__35360\,
            in2 => \_gnd_net_\,
            in3 => \N__35346\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_12\,
            clk => \N__52367\,
            ce => \N__35579\,
            sr => \N__52038\
        );

    \phase_controller_inst1.stoper_tr.counter_13_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35727\,
            in1 => \N__35342\,
            in2 => \_gnd_net_\,
            in3 => \N__35328\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_13\,
            clk => \N__52367\,
            ce => \N__35579\,
            sr => \N__52038\
        );

    \phase_controller_inst1.stoper_tr.counter_14_LC_12_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35711\,
            in1 => \N__35324\,
            in2 => \_gnd_net_\,
            in3 => \N__35310\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_14\,
            clk => \N__52367\,
            ce => \N__35579\,
            sr => \N__52038\
        );

    \phase_controller_inst1.stoper_tr.counter_15_LC_12_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35728\,
            in1 => \N__35561\,
            in2 => \_gnd_net_\,
            in3 => \N__35547\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_15\,
            clk => \N__52367\,
            ce => \N__35579\,
            sr => \N__52038\
        );

    \phase_controller_inst1.stoper_tr.counter_16_LC_12_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35713\,
            in1 => \N__37867\,
            in2 => \_gnd_net_\,
            in3 => \N__35544\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_12_29_0_\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_16\,
            clk => \N__52366\,
            ce => \N__35578\,
            sr => \N__52043\
        );

    \phase_controller_inst1.stoper_tr.counter_17_LC_12_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35717\,
            in1 => \N__37921\,
            in2 => \_gnd_net_\,
            in3 => \N__35541\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_17\,
            clk => \N__52366\,
            ce => \N__35578\,
            sr => \N__52043\
        );

    \phase_controller_inst1.stoper_tr.counter_18_LC_12_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35714\,
            in1 => \N__38343\,
            in2 => \_gnd_net_\,
            in3 => \N__35538\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_18\,
            clk => \N__52366\,
            ce => \N__35578\,
            sr => \N__52043\
        );

    \phase_controller_inst1.stoper_tr.counter_19_LC_12_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35718\,
            in1 => \N__38300\,
            in2 => \_gnd_net_\,
            in3 => \N__35535\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_19\,
            clk => \N__52366\,
            ce => \N__35578\,
            sr => \N__52043\
        );

    \phase_controller_inst1.stoper_tr.counter_20_LC_12_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35715\,
            in1 => \N__35532\,
            in2 => \_gnd_net_\,
            in3 => \N__35514\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_20\,
            clk => \N__52366\,
            ce => \N__35578\,
            sr => \N__52043\
        );

    \phase_controller_inst1.stoper_tr.counter_21_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35719\,
            in1 => \N__35510\,
            in2 => \_gnd_net_\,
            in3 => \N__35490\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_21\,
            clk => \N__52366\,
            ce => \N__35578\,
            sr => \N__52043\
        );

    \phase_controller_inst1.stoper_tr.counter_22_LC_12_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35716\,
            in1 => \N__35487\,
            in2 => \_gnd_net_\,
            in3 => \N__35472\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_22\,
            clk => \N__52366\,
            ce => \N__35578\,
            sr => \N__52043\
        );

    \phase_controller_inst1.stoper_tr.counter_23_LC_12_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35720\,
            in1 => \N__35940\,
            in2 => \_gnd_net_\,
            in3 => \N__35925\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_23\,
            clk => \N__52366\,
            ce => \N__35578\,
            sr => \N__52043\
        );

    \phase_controller_inst1.stoper_tr.counter_24_LC_12_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35721\,
            in1 => \N__35922\,
            in2 => \_gnd_net_\,
            in3 => \N__35904\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_12_30_0_\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_24\,
            clk => \N__52365\,
            ce => \N__35577\,
            sr => \N__52045\
        );

    \phase_controller_inst1.stoper_tr.counter_25_LC_12_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35730\,
            in1 => \N__35900\,
            in2 => \_gnd_net_\,
            in3 => \N__35880\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_25\,
            clk => \N__52365\,
            ce => \N__35577\,
            sr => \N__52045\
        );

    \phase_controller_inst1.stoper_tr.counter_26_LC_12_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35722\,
            in1 => \N__35863\,
            in2 => \_gnd_net_\,
            in3 => \N__35847\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_26\,
            clk => \N__52365\,
            ce => \N__35577\,
            sr => \N__52045\
        );

    \phase_controller_inst1.stoper_tr.counter_27_LC_12_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35731\,
            in1 => \N__35839\,
            in2 => \_gnd_net_\,
            in3 => \N__35817\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_27\,
            clk => \N__52365\,
            ce => \N__35577\,
            sr => \N__52045\
        );

    \phase_controller_inst1.stoper_tr.counter_28_LC_12_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35723\,
            in1 => \N__35806\,
            in2 => \_gnd_net_\,
            in3 => \N__35790\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_28\,
            clk => \N__52365\,
            ce => \N__35577\,
            sr => \N__52045\
        );

    \phase_controller_inst1.stoper_tr.counter_29_LC_12_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35732\,
            in1 => \N__35782\,
            in2 => \_gnd_net_\,
            in3 => \N__35760\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_29\,
            clk => \N__52365\,
            ce => \N__35577\,
            sr => \N__52045\
        );

    \phase_controller_inst1.stoper_tr.counter_30_LC_12_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35724\,
            in1 => \N__35757\,
            in2 => \_gnd_net_\,
            in3 => \N__35739\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_29\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_30\,
            clk => \N__52365\,
            ce => \N__35577\,
            sr => \N__52045\
        );

    \phase_controller_inst1.stoper_tr.counter_31_LC_12_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__35598\,
            in1 => \N__35725\,
            in2 => \_gnd_net_\,
            in3 => \N__35601\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52365\,
            ce => \N__35577\,
            sr => \N__52045\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38213\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.counter_0_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36193\,
            in1 => \N__38151\,
            in2 => \N__38169\,
            in3 => \N__38165\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_0\,
            clk => \N__52467\,
            ce => \N__36058\,
            sr => \N__51928\
        );

    \phase_controller_inst2.stoper_hc.counter_1_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36225\,
            in1 => \N__38133\,
            in2 => \_gnd_net_\,
            in3 => \N__35961\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_1\,
            clk => \N__52467\,
            ce => \N__36058\,
            sr => \N__51928\
        );

    \phase_controller_inst2.stoper_hc.counter_2_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36194\,
            in1 => \N__38604\,
            in2 => \_gnd_net_\,
            in3 => \N__35958\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_2\,
            clk => \N__52467\,
            ce => \N__36058\,
            sr => \N__51928\
        );

    \phase_controller_inst2.stoper_hc.counter_3_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36226\,
            in1 => \N__38586\,
            in2 => \_gnd_net_\,
            in3 => \N__35955\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_3\,
            clk => \N__52467\,
            ce => \N__36058\,
            sr => \N__51928\
        );

    \phase_controller_inst2.stoper_hc.counter_4_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36195\,
            in1 => \N__38568\,
            in2 => \_gnd_net_\,
            in3 => \N__35952\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_4\,
            clk => \N__52467\,
            ce => \N__36058\,
            sr => \N__51928\
        );

    \phase_controller_inst2.stoper_hc.counter_5_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36227\,
            in1 => \N__38550\,
            in2 => \_gnd_net_\,
            in3 => \N__35949\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_5\,
            clk => \N__52467\,
            ce => \N__36058\,
            sr => \N__51928\
        );

    \phase_controller_inst2.stoper_hc.counter_6_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36196\,
            in1 => \N__38529\,
            in2 => \_gnd_net_\,
            in3 => \N__35946\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_6\,
            clk => \N__52467\,
            ce => \N__36058\,
            sr => \N__51928\
        );

    \phase_controller_inst2.stoper_hc.counter_7_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36228\,
            in1 => \N__38505\,
            in2 => \_gnd_net_\,
            in3 => \N__35943\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_7\,
            clk => \N__52467\,
            ce => \N__36058\,
            sr => \N__51928\
        );

    \phase_controller_inst2.stoper_hc.counter_8_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36205\,
            in1 => \N__38484\,
            in2 => \_gnd_net_\,
            in3 => \N__35988\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_8\,
            clk => \N__52462\,
            ce => \N__36076\,
            sr => \N__51933\
        );

    \phase_controller_inst2.stoper_hc.counter_9_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36224\,
            in1 => \N__38463\,
            in2 => \_gnd_net_\,
            in3 => \N__35985\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_9\,
            clk => \N__52462\,
            ce => \N__36076\,
            sr => \N__51933\
        );

    \phase_controller_inst2.stoper_hc.counter_10_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36202\,
            in1 => \N__38733\,
            in2 => \_gnd_net_\,
            in3 => \N__35982\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_10\,
            clk => \N__52462\,
            ce => \N__36076\,
            sr => \N__51933\
        );

    \phase_controller_inst2.stoper_hc.counter_11_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36221\,
            in1 => \N__38712\,
            in2 => \_gnd_net_\,
            in3 => \N__35979\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_11\,
            clk => \N__52462\,
            ce => \N__36076\,
            sr => \N__51933\
        );

    \phase_controller_inst2.stoper_hc.counter_12_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36203\,
            in1 => \N__38691\,
            in2 => \_gnd_net_\,
            in3 => \N__35976\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_12\,
            clk => \N__52462\,
            ce => \N__36076\,
            sr => \N__51933\
        );

    \phase_controller_inst2.stoper_hc.counter_13_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36222\,
            in1 => \N__38667\,
            in2 => \_gnd_net_\,
            in3 => \N__35973\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_13\,
            clk => \N__52462\,
            ce => \N__36076\,
            sr => \N__51933\
        );

    \phase_controller_inst2.stoper_hc.counter_14_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36204\,
            in1 => \N__38646\,
            in2 => \_gnd_net_\,
            in3 => \N__35970\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_14\,
            clk => \N__52462\,
            ce => \N__36076\,
            sr => \N__51933\
        );

    \phase_controller_inst2.stoper_hc.counter_15_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36223\,
            in1 => \N__38625\,
            in2 => \_gnd_net_\,
            in3 => \N__35967\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_15\,
            clk => \N__52462\,
            ce => \N__36076\,
            sr => \N__51933\
        );

    \phase_controller_inst2.stoper_hc.counter_16_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36206\,
            in1 => \N__49957\,
            in2 => \_gnd_net_\,
            in3 => \N__35964\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_16\,
            clk => \N__52458\,
            ce => \N__36077\,
            sr => \N__51934\
        );

    \phase_controller_inst2.stoper_hc.counter_17_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36210\,
            in1 => \N__49981\,
            in2 => \_gnd_net_\,
            in3 => \N__36015\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_17\,
            clk => \N__52458\,
            ce => \N__36077\,
            sr => \N__51934\
        );

    \phase_controller_inst2.stoper_hc.counter_18_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36207\,
            in1 => \N__49843\,
            in2 => \_gnd_net_\,
            in3 => \N__36012\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_18\,
            clk => \N__52458\,
            ce => \N__36077\,
            sr => \N__51934\
        );

    \phase_controller_inst2.stoper_hc.counter_19_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36211\,
            in1 => \N__49865\,
            in2 => \_gnd_net_\,
            in3 => \N__36009\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_19\,
            clk => \N__52458\,
            ce => \N__36077\,
            sr => \N__51934\
        );

    \phase_controller_inst2.stoper_hc.counter_20_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36208\,
            in1 => \N__41288\,
            in2 => \_gnd_net_\,
            in3 => \N__36006\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_20\,
            clk => \N__52458\,
            ce => \N__36077\,
            sr => \N__51934\
        );

    \phase_controller_inst2.stoper_hc.counter_21_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36212\,
            in1 => \N__41315\,
            in2 => \_gnd_net_\,
            in3 => \N__36003\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_21\,
            clk => \N__52458\,
            ce => \N__36077\,
            sr => \N__51934\
        );

    \phase_controller_inst2.stoper_hc.counter_22_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36209\,
            in1 => \N__41642\,
            in2 => \_gnd_net_\,
            in3 => \N__36000\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_22\,
            clk => \N__52458\,
            ce => \N__36077\,
            sr => \N__51934\
        );

    \phase_controller_inst2.stoper_hc.counter_23_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36213\,
            in1 => \N__41678\,
            in2 => \_gnd_net_\,
            in3 => \N__35997\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_23\,
            clk => \N__52458\,
            ce => \N__36077\,
            sr => \N__51934\
        );

    \phase_controller_inst2.stoper_hc.counter_24_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36197\,
            in1 => \N__49771\,
            in2 => \_gnd_net_\,
            in3 => \N__35994\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_24\,
            clk => \N__52452\,
            ce => \N__36084\,
            sr => \N__51940\
        );

    \phase_controller_inst2.stoper_hc.counter_25_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36229\,
            in1 => \N__49789\,
            in2 => \_gnd_net_\,
            in3 => \N__35991\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_25\,
            clk => \N__52452\,
            ce => \N__36084\,
            sr => \N__51940\
        );

    \phase_controller_inst2.stoper_hc.counter_26_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36198\,
            in1 => \N__50305\,
            in2 => \_gnd_net_\,
            in3 => \N__36261\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_26\,
            clk => \N__52452\,
            ce => \N__36084\,
            sr => \N__51940\
        );

    \phase_controller_inst2.stoper_hc.counter_27_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36230\,
            in1 => \N__50276\,
            in2 => \_gnd_net_\,
            in3 => \N__36258\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_27\,
            clk => \N__52452\,
            ce => \N__36084\,
            sr => \N__51940\
        );

    \phase_controller_inst2.stoper_hc.counter_28_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36199\,
            in1 => \N__38934\,
            in2 => \_gnd_net_\,
            in3 => \N__36255\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_28\,
            clk => \N__52452\,
            ce => \N__36084\,
            sr => \N__51940\
        );

    \phase_controller_inst2.stoper_hc.counter_29_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36231\,
            in1 => \N__38898\,
            in2 => \_gnd_net_\,
            in3 => \N__36252\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_29\,
            clk => \N__52452\,
            ce => \N__36084\,
            sr => \N__51940\
        );

    \phase_controller_inst2.stoper_hc.counter_30_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36200\,
            in1 => \N__36249\,
            in2 => \_gnd_net_\,
            in3 => \N__36234\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_29\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_30\,
            clk => \N__52452\,
            ce => \N__36084\,
            sr => \N__51940\
        );

    \phase_controller_inst2.stoper_hc.counter_31_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__36099\,
            in1 => \N__36201\,
            in2 => \_gnd_net_\,
            in3 => \N__36102\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52452\,
            ce => \N__36084\,
            sr => \N__51940\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_28_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47667\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52445\,
            ce => \N__50155\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_22_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37632\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52439\,
            ce => \N__36335\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_26_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37785\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52439\,
            ce => \N__36335\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_15_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37419\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52439\,
            ce => \N__36335\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_27_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37764\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52439\,
            ce => \N__36335\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_20_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37677\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52439\,
            ce => \N__36335\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_23_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37611\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52434\,
            ce => \N__36339\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_7_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37176\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52434\,
            ce => \N__36339\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_18_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37698\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52434\,
            ce => \N__36339\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_16_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37398\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52434\,
            ce => \N__36339\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_19_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__38442\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52434\,
            ce => \N__36339\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_21_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37653\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52434\,
            ce => \N__36339\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_2_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__36653\,
            in1 => \N__36754\,
            in2 => \N__41218\,
            in3 => \N__36795\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52429\,
            ce => 'H',
            sr => \N__51954\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__39157\,
            in1 => \N__39881\,
            in2 => \_gnd_net_\,
            in3 => \N__39909\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001101"
        )
    port map (
            in0 => \N__39908\,
            in1 => \N__39156\,
            in2 => \N__39885\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__39704\,
            in1 => \N__39857\,
            in2 => \_gnd_net_\,
            in3 => \N__39158\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_28_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47660\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52422\,
            ce => \N__43467\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__37738\,
            in1 => \N__36843\,
            in2 => \_gnd_net_\,
            in3 => \N__36821\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52417\,
            ce => 'H',
            sr => \N__51963\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36728\,
            in2 => \_gnd_net_\,
            in3 => \N__36707\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52417\,
            ce => 'H',
            sr => \N__51963\
        );

    \phase_controller_inst1.state_RNO_0_3_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010111001111"
        )
    port map (
            in0 => \N__37102\,
            in1 => \N__36657\,
            in2 => \N__41211\,
            in3 => \N__37091\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.state_ns_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_3_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111110001111"
        )
    port map (
            in0 => \N__36604\,
            in1 => \N__36534\,
            in2 => \N__36516\,
            in3 => \N__36513\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52411\,
            ce => 'H',
            sr => \N__51966\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__37122\,
            in1 => \N__37106\,
            in2 => \N__36881\,
            in3 => \N__36911\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52411\,
            ce => 'H',
            sr => \N__51966\
        );

    \phase_controller_inst1.state_0_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__37082\,
            in1 => \N__38260\,
            in2 => \N__37107\,
            in3 => \N__37092\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52411\,
            ce => 'H',
            sr => \N__51966\
        );

    \phase_controller_inst1.start_timer_tr_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__38261\,
            in1 => \N__37032\,
            in2 => \N__37083\,
            in3 => \N__37047\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52411\,
            ce => 'H',
            sr => \N__51966\
        );

    \phase_controller_inst1.stoper_tr.running_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000101110"
        )
    port map (
            in0 => \N__36877\,
            in1 => \N__37031\,
            in2 => \N__36978\,
            in3 => \N__36912\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52411\,
            ce => 'H',
            sr => \N__51966\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44154\,
            in1 => \N__43953\,
            in2 => \N__44205\,
            in3 => \N__43932\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44177\,
            in1 => \N__44228\,
            in2 => \N__36858\,
            in3 => \N__36855\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__37740\,
            in1 => \_gnd_net_\,
            in2 => \N__36849\,
            in3 => \N__36822\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_158_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39210\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36801\,
            in2 => \N__39604\,
            in3 => \N__42295\,
            lcout => \phase_controller_inst1.stoper_tr.measured_delay_tr_i_31\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__39579\,
            in1 => \N__39578\,
            in2 => \N__46684\,
            in3 => \N__37326\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_1,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40050\,
            in1 => \N__40049\,
            in2 => \N__46688\,
            in3 => \N__37296\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_2,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40035\,
            in1 => \N__40034\,
            in2 => \N__46685\,
            in3 => \N__37266\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_3,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40020\,
            in1 => \N__40019\,
            in2 => \N__46689\,
            in3 => \N__37236\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_4,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40005\,
            in1 => \N__40004\,
            in2 => \N__46686\,
            in3 => \N__37206\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_5,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__39978\,
            in1 => \N__39977\,
            in2 => \N__46690\,
            in3 => \N__37179\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_6,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__39957\,
            in1 => \N__39956\,
            in2 => \N__46687\,
            in3 => \N__37155\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_7,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__39939\,
            in1 => \N__39938\,
            in2 => \N__46842\,
            in3 => \N__37125\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_8,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__39924\,
            in1 => \N__39923\,
            in2 => \N__46839\,
            in3 => \N__37527\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_9,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40200\,
            in1 => \N__40199\,
            in2 => \N__46843\,
            in3 => \N__37506\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_10,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40185\,
            in1 => \N__40184\,
            in2 => \N__46836\,
            in3 => \N__37485\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_11,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40170\,
            in1 => \N__40169\,
            in2 => \N__46840\,
            in3 => \N__37464\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_12,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40155\,
            in1 => \N__40154\,
            in2 => \N__46837\,
            in3 => \N__37443\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_13,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40140\,
            in1 => \N__40139\,
            in2 => \N__46841\,
            in3 => \N__37422\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_14,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40119\,
            in1 => \N__40118\,
            in2 => \N__46838\,
            in3 => \N__37401\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_15,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40101\,
            in1 => \N__40100\,
            in2 => \N__46844\,
            in3 => \N__37380\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_16,
            ltout => OPEN,
            carryin => \bfn_13_21_0_\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40082\,
            in1 => \N__40086\,
            in2 => \N__46872\,
            in3 => \N__37356\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_17,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40065\,
            in1 => \N__40064\,
            in2 => \N__46845\,
            in3 => \N__37683\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_18,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40329\,
            in1 => \N__40328\,
            in2 => \N__46873\,
            in3 => \N__37680\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_19,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40314\,
            in1 => \N__40313\,
            in2 => \N__46846\,
            in3 => \N__37656\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_20,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40299\,
            in1 => \N__40298\,
            in2 => \N__46874\,
            in3 => \N__37635\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_21,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40284\,
            in1 => \N__40283\,
            in2 => \N__46847\,
            in3 => \N__37614\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_22,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40263\,
            in1 => \N__40262\,
            in2 => \N__46875\,
            in3 => \N__37593\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_23,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40245\,
            in1 => \N__40244\,
            in2 => \N__46876\,
            in3 => \N__37572\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_24,
            ltout => OPEN,
            carryin => \bfn_13_22_0_\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40230\,
            in1 => \N__40229\,
            in2 => \N__46878\,
            in3 => \N__37551\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_25,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40215\,
            in1 => \N__40214\,
            in2 => \N__46877\,
            in3 => \N__37767\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_26,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40494\,
            in1 => \N__40493\,
            in2 => \N__46879\,
            in3 => \N__37746\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_27,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37743\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37739\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38054\,
            in1 => \N__42223\,
            in2 => \_gnd_net_\,
            in3 => \N__37713\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__52385\,
            ce => \N__37972\,
            sr => \N__51999\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38088\,
            in1 => \N__42175\,
            in2 => \_gnd_net_\,
            in3 => \N__37710\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__52385\,
            ce => \N__37972\,
            sr => \N__51999\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38055\,
            in1 => \N__40443\,
            in2 => \_gnd_net_\,
            in3 => \N__37707\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__52385\,
            ce => \N__37972\,
            sr => \N__51999\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38089\,
            in1 => \N__40421\,
            in2 => \_gnd_net_\,
            in3 => \N__37704\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__52385\,
            ce => \N__37972\,
            sr => \N__51999\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38056\,
            in1 => \N__40399\,
            in2 => \_gnd_net_\,
            in3 => \N__37701\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__52385\,
            ce => \N__37972\,
            sr => \N__51999\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38090\,
            in1 => \N__40373\,
            in2 => \_gnd_net_\,
            in3 => \N__37812\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__52385\,
            ce => \N__37972\,
            sr => \N__51999\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38057\,
            in1 => \N__40349\,
            in2 => \_gnd_net_\,
            in3 => \N__37809\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__52385\,
            ce => \N__37972\,
            sr => \N__51999\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38091\,
            in1 => \N__40679\,
            in2 => \_gnd_net_\,
            in3 => \N__37806\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__52385\,
            ce => \N__37972\,
            sr => \N__51999\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38075\,
            in1 => \N__40655\,
            in2 => \_gnd_net_\,
            in3 => \N__37803\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__52381\,
            ce => \N__37968\,
            sr => \N__52005\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38087\,
            in1 => \N__40634\,
            in2 => \_gnd_net_\,
            in3 => \N__37800\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__52381\,
            ce => \N__37968\,
            sr => \N__52005\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38072\,
            in1 => \N__40610\,
            in2 => \_gnd_net_\,
            in3 => \N__37797\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__52381\,
            ce => \N__37968\,
            sr => \N__52005\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38084\,
            in1 => \N__40588\,
            in2 => \_gnd_net_\,
            in3 => \N__37794\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__52381\,
            ce => \N__37968\,
            sr => \N__52005\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38073\,
            in1 => \N__40562\,
            in2 => \_gnd_net_\,
            in3 => \N__37791\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__52381\,
            ce => \N__37968\,
            sr => \N__52005\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38085\,
            in1 => \N__40538\,
            in2 => \_gnd_net_\,
            in3 => \N__37788\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__52381\,
            ce => \N__37968\,
            sr => \N__52005\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38074\,
            in1 => \N__40514\,
            in2 => \_gnd_net_\,
            in3 => \N__37839\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__52381\,
            ce => \N__37968\,
            sr => \N__52005\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38086\,
            in1 => \N__40865\,
            in2 => \_gnd_net_\,
            in3 => \N__37836\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__52381\,
            ce => \N__37968\,
            sr => \N__52005\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38076\,
            in1 => \N__40841\,
            in2 => \_gnd_net_\,
            in3 => \N__37833\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_25_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__52377\,
            ce => \N__37973\,
            sr => \N__52012\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38080\,
            in1 => \N__40817\,
            in2 => \_gnd_net_\,
            in3 => \N__37830\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__52377\,
            ce => \N__37973\,
            sr => \N__52012\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38077\,
            in1 => \N__40797\,
            in2 => \_gnd_net_\,
            in3 => \N__37827\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__52377\,
            ce => \N__37973\,
            sr => \N__52012\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38081\,
            in1 => \N__40775\,
            in2 => \_gnd_net_\,
            in3 => \N__37824\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__52377\,
            ce => \N__37973\,
            sr => \N__52012\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38078\,
            in1 => \N__40753\,
            in2 => \_gnd_net_\,
            in3 => \N__37821\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__52377\,
            ce => \N__37973\,
            sr => \N__52012\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38082\,
            in1 => \N__40727\,
            in2 => \_gnd_net_\,
            in3 => \N__37818\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__52377\,
            ce => \N__37973\,
            sr => \N__52012\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38079\,
            in1 => \N__40703\,
            in2 => \_gnd_net_\,
            in3 => \N__37815\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__52377\,
            ce => \N__37973\,
            sr => \N__52012\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38083\,
            in1 => \N__41069\,
            in2 => \_gnd_net_\,
            in3 => \N__38115\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__52377\,
            ce => \N__37973\,
            sr => \N__52012\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38092\,
            in1 => \N__41045\,
            in2 => \_gnd_net_\,
            in3 => \N__38112\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_13_26_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__52374\,
            ce => \N__37974\,
            sr => \N__52021\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38096\,
            in1 => \N__41024\,
            in2 => \_gnd_net_\,
            in3 => \N__38109\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__52374\,
            ce => \N__37974\,
            sr => \N__52021\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38093\,
            in1 => \N__40988\,
            in2 => \_gnd_net_\,
            in3 => \N__38106\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__52374\,
            ce => \N__37974\,
            sr => \N__52021\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38097\,
            in1 => \N__40954\,
            in2 => \_gnd_net_\,
            in3 => \N__38103\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__52374\,
            ce => \N__37974\,
            sr => \N__52021\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38094\,
            in1 => \N__41004\,
            in2 => \_gnd_net_\,
            in3 => \N__38100\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__52374\,
            ce => \N__37974\,
            sr => \N__52021\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__40968\,
            in1 => \N__38095\,
            in2 => \_gnd_net_\,
            in3 => \N__37977\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52374\,
            ce => \N__37974\,
            sr => \N__52021\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011010100"
        )
    port map (
            in0 => \N__37923\,
            in1 => \N__37905\,
            in2 => \N__37890\,
            in3 => \N__37869\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011110101"
        )
    port map (
            in0 => \N__37922\,
            in1 => \N__37904\,
            in2 => \N__37889\,
            in3 => \N__37868\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_19_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38441\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52372\,
            ce => \N__38424\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__38327\,
            in1 => \N__38312\,
            in2 => \N__38301\,
            in3 => \N__38341\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_13_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__38342\,
            in1 => \N__38328\,
            in2 => \N__38313\,
            in3 => \N__38299\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38271\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52368\,
            ce => 'H',
            sr => \N__52039\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40914\,
            in2 => \_gnd_net_\,
            in3 => \N__40887\,
            lcout => \current_shift_inst.timer_s1.N_153_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38219\,
            in2 => \_gnd_net_\,
            in3 => \N__38762\,
            lcout => \phase_controller_inst2.stoper_hc.counter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38139\,
            in2 => \N__41148\,
            in3 => \N__38150\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38121\,
            in2 => \N__41121\,
            in3 => \N__38132\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38592\,
            in2 => \N__41112\,
            in3 => \N__38603\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38574\,
            in2 => \N__41139\,
            in3 => \N__38585\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38556\,
            in2 => \N__41130\,
            in3 => \N__38567\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43245\,
            in2 => \N__38538\,
            in3 => \N__38549\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41103\,
            in2 => \N__38517\,
            in3 => \N__38528\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43236\,
            in2 => \N__38493\,
            in3 => \N__38504\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43383\,
            in2 => \N__38472\,
            in3 => \N__38483\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43200\,
            in2 => \N__38451\,
            in3 => \N__38462\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43227\,
            in2 => \N__38721\,
            in3 => \N__38732\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43269\,
            in2 => \N__38700\,
            in3 => \N__38711\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38690\,
            in1 => \N__43209\,
            in2 => \N__38679\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43392\,
            in2 => \N__38655\,
            in3 => \N__38666\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43257\,
            in2 => \N__38634\,
            in3 => \N__38645\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43218\,
            in2 => \N__38613\,
            in3 => \N__38624\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50004\,
            in2 => \N__49938\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49818\,
            in2 => \N__49896\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41274\,
            in2 => \N__41343\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41259\,
            in2 => \N__41628\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49755\,
            in2 => \N__49806\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49746\,
            in2 => \N__50262\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38883\,
            in2 => \N__38745\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38796\,
            in2 => \N__38787\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38775\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__38896\,
            in1 => \N__38918\,
            in2 => \_gnd_net_\,
            in3 => \N__38932\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__41612\,
            in1 => \N__43500\,
            in2 => \N__41583\,
            in3 => \N__43485\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__38933\,
            in1 => \_gnd_net_\,
            in2 => \N__38919\,
            in3 => \N__38897\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39087\,
            in1 => \N__38877\,
            in2 => \N__38862\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41373\,
            in2 => \N__38853\,
            in3 => \N__39072\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41352\,
            in2 => \N__38844\,
            in3 => \N__39378\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43374\,
            in2 => \N__38835\,
            in3 => \N__39360\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43551\,
            in2 => \N__38826\,
            in3 => \N__39342\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39324\,
            in1 => \N__43350\,
            in2 => \N__38814\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39306\,
            in1 => \N__41097\,
            in2 => \N__38805\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39288\,
            in1 => \N__43515\,
            in2 => \N__39012\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41085\,
            in2 => \N__39003\,
            in3 => \N__39270\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43296\,
            in2 => \N__38994\,
            in3 => \N__39252\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43284\,
            in2 => \N__38985\,
            in3 => \N__39498\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41364\,
            in2 => \N__38976\,
            in3 => \N__39480\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39462\,
            in1 => \N__41385\,
            in2 => \N__38964\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39441\,
            in1 => \N__43338\,
            in2 => \N__38952\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39423\,
            in1 => \N__43326\,
            in2 => \N__38943\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39405\,
            in1 => \N__43362\,
            in2 => \N__39054\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41838\,
            in2 => \N__41784\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41766\,
            in2 => \N__41703\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41535\,
            in2 => \N__41466\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41454\,
            in2 => \N__41859\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39045\,
            in2 => \N__41550\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39120\,
            in2 => \N__39129\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39036\,
            in2 => \N__39030\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39018\,
            in2 => \N__39138\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39234\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO\,
            ltout => \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39213\,
            in3 => \N__39208\,
            lcout => \phase_controller_inst1.stoper_hc.counter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__39705\,
            in1 => \N__39858\,
            in2 => \_gnd_net_\,
            in3 => \N__39159\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011011100"
        )
    port map (
            in0 => \N__39543\,
            in1 => \N__43313\,
            in2 => \N__43578\,
            in3 => \N__39522\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011110101"
        )
    port map (
            in0 => \N__39521\,
            in1 => \N__43574\,
            in2 => \N__43314\,
            in3 => \N__39542\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44097\,
            in1 => \N__39114\,
            in2 => \_gnd_net_\,
            in3 => \N__42744\,
            lcout => \elapsed_time_ns_1_RNILK91B_0_9\,
            ltout => \elapsed_time_ns_1_RNILK91B_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39108\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.counter_0_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39824\,
            in1 => \N__39086\,
            in2 => \N__39104\,
            in3 => \N__39105\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_0\,
            clk => \N__52423\,
            ce => \N__39675\,
            sr => \N__51958\
        );

    \phase_controller_inst1.stoper_hc.counter_1_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39828\,
            in1 => \N__39071\,
            in2 => \_gnd_net_\,
            in3 => \N__39057\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_1\,
            clk => \N__52423\,
            ce => \N__39675\,
            sr => \N__51958\
        );

    \phase_controller_inst1.stoper_hc.counter_2_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39825\,
            in1 => \N__39377\,
            in2 => \_gnd_net_\,
            in3 => \N__39363\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_2\,
            clk => \N__52423\,
            ce => \N__39675\,
            sr => \N__51958\
        );

    \phase_controller_inst1.stoper_hc.counter_3_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39829\,
            in1 => \N__39359\,
            in2 => \_gnd_net_\,
            in3 => \N__39345\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_3\,
            clk => \N__52423\,
            ce => \N__39675\,
            sr => \N__51958\
        );

    \phase_controller_inst1.stoper_hc.counter_4_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39826\,
            in1 => \N__39341\,
            in2 => \_gnd_net_\,
            in3 => \N__39327\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_4\,
            clk => \N__52423\,
            ce => \N__39675\,
            sr => \N__51958\
        );

    \phase_controller_inst1.stoper_hc.counter_5_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39830\,
            in1 => \N__39323\,
            in2 => \_gnd_net_\,
            in3 => \N__39309\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_5\,
            clk => \N__52423\,
            ce => \N__39675\,
            sr => \N__51958\
        );

    \phase_controller_inst1.stoper_hc.counter_6_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39827\,
            in1 => \N__39305\,
            in2 => \_gnd_net_\,
            in3 => \N__39291\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_6\,
            clk => \N__52423\,
            ce => \N__39675\,
            sr => \N__51958\
        );

    \phase_controller_inst1.stoper_hc.counter_7_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39831\,
            in1 => \N__39287\,
            in2 => \_gnd_net_\,
            in3 => \N__39273\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_7\,
            clk => \N__52423\,
            ce => \N__39675\,
            sr => \N__51958\
        );

    \phase_controller_inst1.stoper_hc.counter_8_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39811\,
            in1 => \N__39269\,
            in2 => \_gnd_net_\,
            in3 => \N__39255\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_8\,
            clk => \N__52418\,
            ce => \N__39681\,
            sr => \N__51964\
        );

    \phase_controller_inst1.stoper_hc.counter_9_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39815\,
            in1 => \N__39251\,
            in2 => \_gnd_net_\,
            in3 => \N__39237\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_9\,
            clk => \N__52418\,
            ce => \N__39681\,
            sr => \N__51964\
        );

    \phase_controller_inst1.stoper_hc.counter_10_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39808\,
            in1 => \N__39497\,
            in2 => \_gnd_net_\,
            in3 => \N__39483\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_10\,
            clk => \N__52418\,
            ce => \N__39681\,
            sr => \N__51964\
        );

    \phase_controller_inst1.stoper_hc.counter_11_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39812\,
            in1 => \N__39479\,
            in2 => \_gnd_net_\,
            in3 => \N__39465\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_11\,
            clk => \N__52418\,
            ce => \N__39681\,
            sr => \N__51964\
        );

    \phase_controller_inst1.stoper_hc.counter_12_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39809\,
            in1 => \N__39458\,
            in2 => \_gnd_net_\,
            in3 => \N__39444\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_12\,
            clk => \N__52418\,
            ce => \N__39681\,
            sr => \N__51964\
        );

    \phase_controller_inst1.stoper_hc.counter_13_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39813\,
            in1 => \N__39440\,
            in2 => \_gnd_net_\,
            in3 => \N__39426\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_13\,
            clk => \N__52418\,
            ce => \N__39681\,
            sr => \N__51964\
        );

    \phase_controller_inst1.stoper_hc.counter_14_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39810\,
            in1 => \N__39422\,
            in2 => \_gnd_net_\,
            in3 => \N__39408\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_14\,
            clk => \N__52418\,
            ce => \N__39681\,
            sr => \N__51964\
        );

    \phase_controller_inst1.stoper_hc.counter_15_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39814\,
            in1 => \N__39404\,
            in2 => \_gnd_net_\,
            in3 => \N__39390\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_15\,
            clk => \N__52418\,
            ce => \N__39681\,
            sr => \N__51964\
        );

    \phase_controller_inst1.stoper_hc.counter_16_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39800\,
            in1 => \N__41798\,
            in2 => \_gnd_net_\,
            in3 => \N__39387\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_16\,
            clk => \N__52412\,
            ce => \N__39679\,
            sr => \N__51967\
        );

    \phase_controller_inst1.stoper_hc.counter_17_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39804\,
            in1 => \N__41825\,
            in2 => \_gnd_net_\,
            in3 => \N__39384\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_17\,
            clk => \N__52412\,
            ce => \N__39679\,
            sr => \N__51967\
        );

    \phase_controller_inst1.stoper_hc.counter_18_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39801\,
            in1 => \N__41717\,
            in2 => \_gnd_net_\,
            in3 => \N__39381\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_18\,
            clk => \N__52412\,
            ce => \N__39679\,
            sr => \N__51967\
        );

    \phase_controller_inst1.stoper_hc.counter_19_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39805\,
            in1 => \N__41744\,
            in2 => \_gnd_net_\,
            in3 => \N__39564\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_19\,
            clk => \N__52412\,
            ce => \N__39679\,
            sr => \N__51967\
        );

    \phase_controller_inst1.stoper_hc.counter_20_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39802\,
            in1 => \N__41480\,
            in2 => \_gnd_net_\,
            in3 => \N__39561\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_20\,
            clk => \N__52412\,
            ce => \N__39679\,
            sr => \N__51967\
        );

    \phase_controller_inst1.stoper_hc.counter_21_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39806\,
            in1 => \N__41501\,
            in2 => \_gnd_net_\,
            in3 => \N__39558\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_21\,
            clk => \N__52412\,
            ce => \N__39679\,
            sr => \N__51967\
        );

    \phase_controller_inst1.stoper_hc.counter_22_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39803\,
            in1 => \N__41399\,
            in2 => \_gnd_net_\,
            in3 => \N__39555\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_22\,
            clk => \N__52412\,
            ce => \N__39679\,
            sr => \N__51967\
        );

    \phase_controller_inst1.stoper_hc.counter_23_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39807\,
            in1 => \N__41426\,
            in2 => \_gnd_net_\,
            in3 => \N__39552\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_23\,
            clk => \N__52412\,
            ce => \N__39679\,
            sr => \N__51967\
        );

    \phase_controller_inst1.stoper_hc.counter_24_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39816\,
            in1 => \N__41564\,
            in2 => \_gnd_net_\,
            in3 => \N__39549\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_24\,
            clk => \N__52407\,
            ce => \N__39680\,
            sr => \N__51973\
        );

    \phase_controller_inst1.stoper_hc.counter_25_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39820\,
            in1 => \N__41605\,
            in2 => \_gnd_net_\,
            in3 => \N__39546\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_25\,
            clk => \N__52407\,
            ce => \N__39680\,
            sr => \N__51973\
        );

    \phase_controller_inst1.stoper_hc.counter_26_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39817\,
            in1 => \N__39541\,
            in2 => \_gnd_net_\,
            in3 => \N__39525\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_26\,
            clk => \N__52407\,
            ce => \N__39680\,
            sr => \N__51973\
        );

    \phase_controller_inst1.stoper_hc.counter_27_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39821\,
            in1 => \N__39515\,
            in2 => \_gnd_net_\,
            in3 => \N__39501\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_27\,
            clk => \N__52407\,
            ce => \N__39680\,
            sr => \N__51973\
        );

    \phase_controller_inst1.stoper_hc.counter_28_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39818\,
            in1 => \N__39902\,
            in2 => \_gnd_net_\,
            in3 => \N__39888\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_28\,
            clk => \N__52407\,
            ce => \N__39680\,
            sr => \N__51973\
        );

    \phase_controller_inst1.stoper_hc.counter_29_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39822\,
            in1 => \N__39875\,
            in2 => \_gnd_net_\,
            in3 => \N__39861\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_29\,
            clk => \N__52407\,
            ce => \N__39680\,
            sr => \N__51973\
        );

    \phase_controller_inst1.stoper_hc.counter_30_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39819\,
            in1 => \N__39850\,
            in2 => \_gnd_net_\,
            in3 => \N__39834\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_29\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_30\,
            clk => \N__52407\,
            ce => \N__39680\,
            sr => \N__51973\
        );

    \phase_controller_inst1.stoper_hc.counter_31_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39823\,
            in1 => \N__39697\,
            in2 => \_gnd_net_\,
            in3 => \N__39708\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52407\,
            ce => \N__39680\,
            sr => \N__51973\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42281\,
            in2 => \N__39630\,
            in3 => \N__42197\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1\,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39621\,
            in2 => \_gnd_net_\,
            in3 => \N__42104\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42366\,
            in2 => \_gnd_net_\,
            in3 => \N__39582\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43830\,
            in2 => \_gnd_net_\,
            in3 => \N__39567\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42447\,
            in3 => \N__40038\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42018\,
            in3 => \N__40023\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42324\,
            in2 => \_gnd_net_\,
            in3 => \N__40008\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42345\,
            in2 => \_gnd_net_\,
            in3 => \N__39993\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39990\,
            in2 => \_gnd_net_\,
            in3 => \N__39960\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0\,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42543\,
            in2 => \_gnd_net_\,
            in3 => \N__39942\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41871\,
            in2 => \_gnd_net_\,
            in3 => \N__39927\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41970\,
            in2 => \_gnd_net_\,
            in3 => \N__39912\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42078\,
            in2 => \_gnd_net_\,
            in3 => \N__40188\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42528\,
            in2 => \_gnd_net_\,
            in3 => \N__40173\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43719\,
            in2 => \_gnd_net_\,
            in3 => \N__40158\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42351\,
            in2 => \_gnd_net_\,
            in3 => \N__40143\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41955\,
            in2 => \_gnd_net_\,
            in3 => \N__40122\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0\,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42474\,
            in2 => \_gnd_net_\,
            in3 => \N__40104\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43140\,
            in2 => \_gnd_net_\,
            in3 => \N__40089\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42429\,
            in2 => \_gnd_net_\,
            in3 => \N__40068\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42057\,
            in2 => \_gnd_net_\,
            in3 => \N__40053\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42597\,
            in2 => \_gnd_net_\,
            in3 => \N__40317\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42582\,
            in2 => \_gnd_net_\,
            in3 => \N__40302\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42468\,
            in2 => \_gnd_net_\,
            in3 => \N__40287\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42453\,
            in2 => \_gnd_net_\,
            in3 => \N__40266\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0\,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41943\,
            in2 => \_gnd_net_\,
            in3 => \N__40248\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42552\,
            in2 => \_gnd_net_\,
            in3 => \N__40233\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42858\,
            in2 => \_gnd_net_\,
            in3 => \N__40218\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42843\,
            in2 => \_gnd_net_\,
            in3 => \N__40203\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42558\,
            in2 => \_gnd_net_\,
            in3 => \N__40482\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__42294\,
            in1 => \N__40479\,
            in2 => \_gnd_net_\,
            in3 => \N__40473\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40441\,
            in2 => \N__42230\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__52386\,
            ce => \N__42147\,
            sr => \N__52000\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40420\,
            in2 => \N__42182\,
            in3 => \N__40446\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__52386\,
            ce => \N__42147\,
            sr => \N__52000\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40442\,
            in2 => \N__40400\,
            in3 => \N__40428\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__52386\,
            ce => \N__42147\,
            sr => \N__52000\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40372\,
            in2 => \N__40425\,
            in3 => \N__40404\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__52386\,
            ce => \N__42147\,
            sr => \N__52000\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40348\,
            in2 => \N__40401\,
            in3 => \N__40380\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__52386\,
            ce => \N__42147\,
            sr => \N__52000\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40678\,
            in2 => \N__40377\,
            in3 => \N__40356\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__52386\,
            ce => \N__42147\,
            sr => \N__52000\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40654\,
            in2 => \N__40353\,
            in3 => \N__40332\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__52386\,
            ce => \N__42147\,
            sr => \N__52000\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40633\,
            in2 => \N__40683\,
            in3 => \N__40662\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__52386\,
            ce => \N__42147\,
            sr => \N__52000\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40609\,
            in2 => \N__40659\,
            in3 => \N__40638\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_14_25_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__52382\,
            ce => \N__42157\,
            sr => \N__52006\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40635\,
            in2 => \N__40589\,
            in3 => \N__40617\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__52382\,
            ce => \N__42157\,
            sr => \N__52006\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40561\,
            in2 => \N__40614\,
            in3 => \N__40593\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__52382\,
            ce => \N__42157\,
            sr => \N__52006\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40537\,
            in2 => \N__40590\,
            in3 => \N__40569\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__52382\,
            ce => \N__42157\,
            sr => \N__52006\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40513\,
            in2 => \N__40566\,
            in3 => \N__40545\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__52382\,
            ce => \N__42157\,
            sr => \N__52006\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40864\,
            in2 => \N__40542\,
            in3 => \N__40521\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__52382\,
            ce => \N__42157\,
            sr => \N__52006\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40840\,
            in2 => \N__40518\,
            in3 => \N__40497\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__52382\,
            ce => \N__42157\,
            sr => \N__52006\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40816\,
            in2 => \N__40869\,
            in3 => \N__40848\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__52382\,
            ce => \N__42157\,
            sr => \N__52006\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40795\,
            in2 => \N__40845\,
            in3 => \N__40824\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_14_26_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__52378\,
            ce => \N__42159\,
            sr => \N__52013\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40774\,
            in2 => \N__40821\,
            in3 => \N__40800\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__52378\,
            ce => \N__42159\,
            sr => \N__52013\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40796\,
            in2 => \N__40754\,
            in3 => \N__40782\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__52378\,
            ce => \N__42159\,
            sr => \N__52013\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40726\,
            in2 => \N__40779\,
            in3 => \N__40758\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__52378\,
            ce => \N__42159\,
            sr => \N__52013\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40702\,
            in2 => \N__40755\,
            in3 => \N__40734\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__52378\,
            ce => \N__42159\,
            sr => \N__52013\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41068\,
            in2 => \N__40731\,
            in3 => \N__40710\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__52378\,
            ce => \N__42159\,
            sr => \N__52013\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41044\,
            in2 => \N__40707\,
            in3 => \N__40686\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__52378\,
            ce => \N__42159\,
            sr => \N__52013\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41023\,
            in2 => \N__41073\,
            in3 => \N__41052\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__52378\,
            ce => \N__42159\,
            sr => \N__52013\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40987\,
            in2 => \N__41049\,
            in3 => \N__41028\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_14_27_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__52375\,
            ce => \N__42158\,
            sr => \N__52022\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41025\,
            in2 => \N__40955\,
            in3 => \N__41007\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__52375\,
            ce => \N__42158\,
            sr => \N__52022\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41003\,
            in2 => \N__40992\,
            in3 => \N__40971\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__52375\,
            ce => \N__42158\,
            sr => \N__52022\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40967\,
            in2 => \N__40956\,
            in3 => \N__40935\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__52375\,
            ce => \N__42158\,
            sr => \N__52022\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40932\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52375\,
            ce => \N__42158\,
            sr => \N__52022\
        );

    \phase_controller_inst1.S1_LC_14_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41229\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52371\,
            ce => 'H',
            sr => \N__52035\
        );

    \current_shift_inst.timer_s1.running_LC_14_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__41169\,
            in1 => \N__40921\,
            in2 => \_gnd_net_\,
            in3 => \N__40892\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52369\,
            ce => 'H',
            sr => \N__52040\
        );

    \current_shift_inst.stop_timer_s1_LC_14_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__41227\,
            in1 => \N__41243\,
            in2 => \N__41172\,
            in3 => \N__40891\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52369\,
            ce => 'H',
            sr => \N__52040\
        );

    \current_shift_inst.start_timer_s1_LC_14_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__41242\,
            in1 => \N__41170\,
            in2 => \_gnd_net_\,
            in3 => \N__41228\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52369\,
            ce => 'H',
            sr => \N__52040\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_0_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47643\,
            in2 => \_gnd_net_\,
            in3 => \N__47149\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52475\,
            ce => \N__50147\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_3_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45722\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52475\,
            ce => \N__50147\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_4_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45701\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52475\,
            ce => \N__50147\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_1_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45764\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52475\,
            ce => \N__50147\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_2_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45743\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52475\,
            ce => \N__50147\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_6_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45935\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52475\,
            ce => \N__50147\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_6_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45939\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52468\,
            ce => \N__43456\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_8_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45900\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52468\,
            ce => \N__43456\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_12_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45834\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52468\,
            ce => \N__43456\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45768\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52468\,
            ce => \N__43456\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_11_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45852\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52468\,
            ce => \N__43456\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_2_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45747\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52468\,
            ce => \N__43456\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__41331\,
            in1 => \N__41322\,
            in2 => \N__41301\,
            in3 => \N__41268\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_20_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45992\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52463\,
            ce => \N__50145\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__41330\,
            in1 => \N__41321\,
            in2 => \N__41300\,
            in3 => \N__41267\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_21_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45975\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52463\,
            ce => \N__50145\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__41685\,
            in1 => \N__41664\,
            in2 => \N__41655\,
            in3 => \N__45789\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_22_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46940\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52463\,
            ce => \N__50145\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__41684\,
            in1 => \N__41663\,
            in2 => \N__41654\,
            in3 => \N__45788\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__41616\,
            in1 => \N__43499\,
            in2 => \N__41582\,
            in3 => \N__43484\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001110"
        )
    port map (
            in0 => \N__43560\,
            in1 => \N__41523\,
            in2 => \N__41513\,
            in3 => \N__41487\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_20_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45996\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52453\,
            ce => \N__43468\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111010101111"
        )
    port map (
            in0 => \N__43559\,
            in1 => \N__41522\,
            in2 => \N__41514\,
            in3 => \N__41486\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__41442\,
            in1 => \N__41433\,
            in2 => \N__41411\,
            in3 => \N__41847\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_22_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46944\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52453\,
            ce => \N__43468\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__41441\,
            in1 => \N__41432\,
            in2 => \N__41412\,
            in3 => \N__41846\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_23_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46923\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52453\,
            ce => \N__43468\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__43539\,
            in1 => \N__41832\,
            in2 => \N__41811\,
            in3 => \N__41775\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__43538\,
            in1 => \N__41831\,
            in2 => \N__41810\,
            in3 => \N__41774\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_17_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49923\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52446\,
            ce => \N__43470\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__41760\,
            in1 => \N__41751\,
            in2 => \N__41730\,
            in3 => \N__43527\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_18_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49578\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52446\,
            ce => \N__43470\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__41759\,
            in1 => \N__41750\,
            in2 => \N__41729\,
            in3 => \N__43526\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50343\,
            in1 => \N__41691\,
            in2 => \_gnd_net_\,
            in3 => \N__50822\,
            lcout => \elapsed_time_ns_1_RNIK63T9_0_8\,
            ltout => \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41910\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41907\,
            in1 => \N__48090\,
            in2 => \_gnd_net_\,
            in3 => \N__50825\,
            lcout => \elapsed_time_ns_1_RNI69DN9_0_28\,
            ltout => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41901\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41898\,
            in1 => \N__47916\,
            in2 => \_gnd_net_\,
            in3 => \N__50824\,
            lcout => \elapsed_time_ns_1_RNIU0DN9_0_20\,
            ltout => \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41892\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41889\,
            in1 => \N__47868\,
            in2 => \_gnd_net_\,
            in3 => \N__50823\,
            lcout => \elapsed_time_ns_1_RNIL73T9_0_9\,
            ltout => \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41883\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41880\,
            in1 => \N__42807\,
            in2 => \_gnd_net_\,
            in3 => \N__44098\,
            lcout => \elapsed_time_ns_1_RNIU7OBB_0_11\,
            ltout => \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41874\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41988\,
            in1 => \N__47937\,
            in2 => \_gnd_net_\,
            in3 => \N__50836\,
            lcout => \elapsed_time_ns_1_RNI68CN9_0_19\,
            ltout => \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41982\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50837\,
            in1 => \N__43659\,
            in2 => \_gnd_net_\,
            in3 => \N__48063\,
            lcout => \elapsed_time_ns_1_RNIV2EN9_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41979\,
            in1 => \N__42768\,
            in2 => \_gnd_net_\,
            in3 => \N__44099\,
            lcout => \elapsed_time_ns_1_RNIV8OBB_0_12\,
            ltout => \elapsed_time_ns_1_RNIV8OBB_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41973\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41930\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42044\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44071\,
            in1 => \N__41931\,
            in2 => \_gnd_net_\,
            in3 => \N__42672\,
            lcout => \elapsed_time_ns_1_RNI4EOBB_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42702\,
            in1 => \N__41919\,
            in2 => \_gnd_net_\,
            in3 => \N__44069\,
            lcout => \elapsed_time_ns_1_RNI0AOBB_0_13\,
            ltout => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41913\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42872\,
            in1 => \N__42918\,
            in2 => \_gnd_net_\,
            in3 => \N__44073\,
            lcout => \elapsed_time_ns_1_RNI6HPBB_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44070\,
            in1 => \N__42066\,
            in2 => \_gnd_net_\,
            in3 => \N__43110\,
            lcout => \elapsed_time_ns_1_RNIV9PBB_0_21\,
            ltout => \elapsed_time_ns_1_RNIV9PBB_0_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42060\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44072\,
            in1 => \N__42045\,
            in2 => \_gnd_net_\,
            in3 => \N__42957\,
            lcout => \elapsed_time_ns_1_RNI4FPBB_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__44264\,
            in1 => \N__42240\,
            in2 => \N__42006\,
            in3 => \N__42819\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__42314\,
            in1 => \N__42681\,
            in2 => \N__42033\,
            in3 => \N__43047\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42027\,
            in2 => \N__42030\,
            in3 => \N__42837\,
            lcout => \elapsed_time_ns_1_RNIIH91B_0_6\,
            ltout => \elapsed_time_ns_1_RNIIH91B_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42021\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42005\,
            in1 => \N__42333\,
            in2 => \_gnd_net_\,
            in3 => \N__44043\,
            lcout => \elapsed_time_ns_1_RNIJI91B_0_7\,
            ltout => \elapsed_time_ns_1_RNIJI91B_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42327\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42280\,
            in1 => \N__42315\,
            in2 => \_gnd_net_\,
            in3 => \N__44044\,
            lcout => \elapsed_time_ns_1_RNI0CQBB_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42092\,
            in1 => \N__42113\,
            in2 => \N__43862\,
            in3 => \N__42206\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42234\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52413\,
            ce => \N__42135\,
            sr => \N__51968\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42198\,
            in1 => \N__42207\,
            in2 => \_gnd_net_\,
            in3 => \N__44092\,
            lcout => \elapsed_time_ns_1_RNIDC91B_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42186\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52413\,
            ce => \N__42135\,
            sr => \N__51968\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42105\,
            in1 => \N__42114\,
            in2 => \_gnd_net_\,
            in3 => \N__44093\,
            lcout => \elapsed_time_ns_1_RNIED91B_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44094\,
            in1 => \N__42378\,
            in2 => \_gnd_net_\,
            in3 => \N__42093\,
            lcout => \elapsed_time_ns_1_RNIFE91B_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44279\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44104\,
            in1 => \N__42438\,
            in2 => \_gnd_net_\,
            in3 => \N__43128\,
            lcout => \elapsed_time_ns_1_RNIU8PBB_0_20\,
            ltout => \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42432\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__42417\,
            in1 => \N__44444\,
            in2 => \_gnd_net_\,
            in3 => \N__44348\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_156_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42377\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44103\,
            in1 => \N__42360\,
            in2 => \_gnd_net_\,
            in3 => \N__42651\,
            lcout => \elapsed_time_ns_1_RNI3DOBB_0_16\,
            ltout => \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42354\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44240\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42339\,
            in1 => \N__42786\,
            in2 => \_gnd_net_\,
            in3 => \N__44100\,
            lcout => \elapsed_time_ns_1_RNIT6OBB_0_10\,
            ltout => \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42546\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44101\,
            in1 => \N__42723\,
            in2 => \_gnd_net_\,
            in3 => \N__42537\,
            lcout => \elapsed_time_ns_1_RNI1BOBB_0_14\,
            ltout => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42531\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42521\,
            in1 => \N__44552\,
            in2 => \N__44510\,
            in3 => \N__42504\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42483\,
            in1 => \N__42630\,
            in2 => \_gnd_net_\,
            in3 => \N__44102\,
            lcout => \elapsed_time_ns_1_RNI5FOBB_0_18\,
            ltout => \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42477\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42575\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__42462\,
            in1 => \N__44109\,
            in2 => \_gnd_net_\,
            in3 => \N__42939\,
            lcout => \elapsed_time_ns_1_RNI3EPBB_0_25\,
            ltout => \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42456\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42606\,
            in1 => \N__43074\,
            in2 => \_gnd_net_\,
            in3 => \N__44107\,
            lcout => \elapsed_time_ns_1_RNI0BPBB_0_22\,
            ltout => \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42600\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42591\,
            in1 => \N__43038\,
            in2 => \_gnd_net_\,
            in3 => \N__44108\,
            lcout => \elapsed_time_ns_1_RNI1CPBB_0_23\,
            ltout => \elapsed_time_ns_1_RNI1CPBB_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42585\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42576\,
            in1 => \N__43002\,
            in2 => \_gnd_net_\,
            in3 => \N__44110\,
            lcout => \elapsed_time_ns_1_RNI2DPBB_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44112\,
            in1 => \N__42567\,
            in2 => \_gnd_net_\,
            in3 => \N__42981\,
            lcout => \elapsed_time_ns_1_RNIVAQBB_0_30\,
            ltout => \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42561\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43968\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__45011\,
            in1 => \N__45406\,
            in2 => \_gnd_net_\,
            in3 => \N__44949\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42876\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42852\,
            in1 => \N__43020\,
            in2 => \_gnd_net_\,
            in3 => \N__44111\,
            lcout => \elapsed_time_ns_1_RNI7IPBB_0_29\,
            ltout => \elapsed_time_ns_1_RNI7IPBB_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42846\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__42830\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44291\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42797\,
            in1 => \N__42779\,
            in2 => \N__42761\,
            in3 => \N__42734\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42716\,
            in2 => \N__42705\,
            in3 => \N__42692\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42662\,
            in1 => \N__42641\,
            in2 => \N__43745\,
            in3 => \N__42623\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42612\,
            in1 => \N__43088\,
            in2 => \_gnd_net_\,
            in3 => \N__44106\,
            lcout => \elapsed_time_ns_1_RNI6GOBB_0_19\,
            ltout => \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43143\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43121\,
            in1 => \N__43100\,
            in2 => \N__43089\,
            in3 => \N__43067\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43056\,
            in1 => \N__42963\,
            in2 => \N__43050\,
            in3 => \N__42897\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43031\,
            in1 => \N__43013\,
            in2 => \N__42998\,
            in3 => \N__42974\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44123\,
            in1 => \N__42950\,
            in2 => \N__42935\,
            in3 => \N__42908\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_15_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__51149\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44711\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_15_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51300\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_28_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_15_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42891\,
            in2 => \_gnd_net_\,
            in3 => \N__42879\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_15_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43191\,
            in2 => \_gnd_net_\,
            in3 => \N__43176\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_15_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43173\,
            in2 => \_gnd_net_\,
            in3 => \N__43161\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_15_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44784\,
            in2 => \_gnd_net_\,
            in3 => \N__43158\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_15_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46829\,
            in2 => \N__45315\,
            in3 => \N__43155\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_15_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45261\,
            in2 => \N__46880\,
            in3 => \N__43152\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_15_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45213\,
            in2 => \N__46881\,
            in3 => \N__43149\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_15_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45174\,
            in2 => \_gnd_net_\,
            in3 => \N__43146\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\,
            ltout => OPEN,
            carryin => \bfn_15_29_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_LC_15_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45132\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_LC_15_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45087\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_LC_15_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45039\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_LC_15_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45642\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_LC_15_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45591\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_LC_15_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45561\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_LC_15_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45531\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_LC_15_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45507\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_30_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_LC_15_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45480\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_LC_15_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45450\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_LC_15_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45363\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_15_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43272\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_11_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45851\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52480\,
            ce => \N__50146\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_14_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46038\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52480\,
            ce => \N__50146\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_5_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45953\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52480\,
            ce => \N__50146\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_7_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45914\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52480\,
            ce => \N__50146\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_10_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45866\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52476\,
            ce => \N__50131\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_15_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46022\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52476\,
            ce => \N__50131\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_12_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45830\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52476\,
            ce => \N__50131\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_9_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45881\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52476\,
            ce => \N__50131\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_13_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46052\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52476\,
            ce => \N__50131\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_8_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45896\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52476\,
            ce => \N__50131\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_3_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45723\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52469\,
            ce => \N__43435\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_15_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46023\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52469\,
            ce => \N__43435\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_5_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45957\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52469\,
            ce => \N__43435\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_13_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46053\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52469\,
            ce => \N__43435\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_14_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46037\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52469\,
            ce => \N__43435\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_27_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50246\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52469\,
            ce => \N__43435\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_9_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45882\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52469\,
            ce => \N__43435\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_10_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45867\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52469\,
            ce => \N__43435\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_26_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50225\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52464\,
            ce => \N__43469\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_21_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45974\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52464\,
            ce => \N__43469\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_4_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45702\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52464\,
            ce => \N__43469\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_16_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49589\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52464\,
            ce => \N__43469\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_19_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50015\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52464\,
            ce => \N__43469\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_7_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45918\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52464\,
            ce => \N__43469\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_24_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50204\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52464\,
            ce => \N__43469\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_25_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50183\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52464\,
            ce => \N__43469\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43674\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43611\,
            in1 => \N__47961\,
            in2 => \_gnd_net_\,
            in3 => \N__50847\,
            lcout => \elapsed_time_ns_1_RNI57CN9_0_18\,
            ltout => \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43605\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50715\,
            in1 => \N__43602\,
            in2 => \_gnd_net_\,
            in3 => \N__50846\,
            lcout => \elapsed_time_ns_1_RNIF13T9_0_3\,
            ltout => \elapsed_time_ns_1_RNIF13T9_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43596\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50325\,
            in1 => \N__43593\,
            in2 => \_gnd_net_\,
            in3 => \N__50850\,
            lcout => \elapsed_time_ns_1_RNIJ53T9_0_7\,
            ltout => \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43587\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46095\,
            in1 => \N__50646\,
            in2 => \_gnd_net_\,
            in3 => \N__50848\,
            lcout => \elapsed_time_ns_1_RNIDV2T9_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50849\,
            in1 => \N__46073\,
            in2 => \_gnd_net_\,
            in3 => \N__50601\,
            lcout => \elapsed_time_ns_1_RNIE03T9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43584\,
            in1 => \N__48000\,
            in2 => \_gnd_net_\,
            in3 => \N__50852\,
            lcout => \elapsed_time_ns_1_RNI35CN9_0_16\,
            ltout => \elapsed_time_ns_1_RNI35CN9_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43647\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43644\,
            in1 => \N__47847\,
            in2 => \_gnd_net_\,
            in3 => \N__50851\,
            lcout => \elapsed_time_ns_1_RNITUBN9_0_10\,
            ltout => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43638\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43703\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50697\,
            in1 => \N__43635\,
            in2 => \_gnd_net_\,
            in3 => \N__50815\,
            lcout => \elapsed_time_ns_1_RNIG23T9_0_4\,
            ltout => \elapsed_time_ns_1_RNIG23T9_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43629\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43626\,
            in1 => \N__48018\,
            in2 => \_gnd_net_\,
            in3 => \N__50817\,
            lcout => \elapsed_time_ns_1_RNI24CN9_0_15\,
            ltout => \elapsed_time_ns_1_RNI24CN9_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43620\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43617\,
            in1 => \N__48039\,
            in2 => \_gnd_net_\,
            in3 => \N__50816\,
            lcout => \elapsed_time_ns_1_RNI13CN9_0_14\,
            ltout => \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43707\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43704\,
            in1 => \N__48144\,
            in2 => \_gnd_net_\,
            in3 => \N__50818\,
            lcout => \elapsed_time_ns_1_RNI25DN9_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43695\,
            in1 => \N__47826\,
            in2 => \_gnd_net_\,
            in3 => \N__50833\,
            lcout => \elapsed_time_ns_1_RNIUVBN9_0_11\,
            ltout => \elapsed_time_ns_1_RNIUVBN9_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43689\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47979\,
            in1 => \N__43686\,
            in2 => \_gnd_net_\,
            in3 => \N__50834\,
            lcout => \elapsed_time_ns_1_RNI46CN9_0_17\,
            ltout => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43680\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43785\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__43758\,
            in1 => \N__50907\,
            in2 => \N__43881\,
            in3 => \N__48326\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__43673\,
            in1 => \_gnd_net_\,
            in2 => \N__43677\,
            in3 => \N__50370\,
            lcout => \elapsed_time_ns_1_RNII43T9_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43658\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43770\,
            in1 => \N__48168\,
            in2 => \_gnd_net_\,
            in3 => \N__50845\,
            lcout => \elapsed_time_ns_1_RNI03DN9_0_22\,
            ltout => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43764\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47822\,
            in1 => \N__47840\,
            in2 => \N__50057\,
            in3 => \N__47861\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48032\,
            in2 => \N__43761\,
            in3 => \N__50426\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43800\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43752\,
            in1 => \N__43728\,
            in2 => \_gnd_net_\,
            in3 => \N__44074\,
            lcout => \elapsed_time_ns_1_RNI2COBB_0_15\,
            ltout => \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43722\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47975\,
            in1 => \N__47993\,
            in2 => \N__47957\,
            in3 => \N__48014\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43811\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47894\,
            in1 => \N__47909\,
            in2 => \N__48167\,
            in3 => \N__47930\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43890\,
            in1 => \N__43869\,
            in2 => \N__43884\,
            in3 => \N__43818\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__50396\,
            in1 => \N__48104\,
            in2 => \N__48123\,
            in3 => \N__48080\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43863\,
            in1 => \N__43839\,
            in2 => \_gnd_net_\,
            in3 => \N__44042\,
            lcout => \elapsed_time_ns_1_RNIGF91B_0_4\,
            ltout => \elapsed_time_ns_1_RNIGF91B_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43833\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__50891\,
            in1 => \N__48137\,
            in2 => \N__48059\,
            in3 => \N__50477\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43812\,
            in1 => \N__48105\,
            in2 => \_gnd_net_\,
            in3 => \N__50873\,
            lcout => \elapsed_time_ns_1_RNI47DN9_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48122\,
            in2 => \N__50880\,
            in3 => \N__43799\,
            lcout => \elapsed_time_ns_1_RNI36DN9_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47895\,
            in1 => \N__43784\,
            in2 => \_gnd_net_\,
            in3 => \N__50869\,
            lcout => \elapsed_time_ns_1_RNIV1DN9_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44448\,
            in2 => \_gnd_net_\,
            in3 => \N__44349\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_155_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44280\,
            in1 => \N__44301\,
            in2 => \_gnd_net_\,
            in3 => \N__44095\,
            lcout => \elapsed_time_ns_1_RNIHG91B_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44241\,
            in1 => \N__44268\,
            in2 => \_gnd_net_\,
            in3 => \N__44096\,
            lcout => \elapsed_time_ns_1_RNIKJ91B_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44229\,
            in1 => \N__44201\,
            in2 => \N__44181\,
            in3 => \N__44153\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43967\,
            in1 => \N__44133\,
            in2 => \_gnd_net_\,
            in3 => \N__44105\,
            lcout => \elapsed_time_ns_1_RNI5GPBB_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44648\,
            in1 => \N__43952\,
            in2 => \N__44604\,
            in3 => \N__43931\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44565\,
            in1 => \N__43911\,
            in2 => \N__44538\,
            in3 => \N__44577\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43905\,
            in1 => \N__43899\,
            in2 => \N__43893\,
            in3 => \N__44355\,
            lcout => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44603\,
            in1 => \N__44409\,
            in2 => \N__44388\,
            in3 => \N__44576\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44564\,
            in2 => \_gnd_net_\,
            in3 => \N__44553\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44528\,
            in2 => \_gnd_net_\,
            in3 => \N__44486\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44529\,
            in1 => \N__44514\,
            in2 => \N__44490\,
            in3 => \N__44475\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44634\,
            in1 => \N__44469\,
            in2 => \N__44463\,
            in3 => \N__44460\,
            lcout => \current_shift_inst.PI_CTRL.N_150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44437\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44402\,
            in2 => \_gnd_net_\,
            in3 => \N__44387\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44687\,
            in1 => \N__44669\,
            in2 => \N__44358\,
            in3 => \N__44699\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44700\,
            in1 => \N__44688\,
            in2 => \N__44673\,
            in3 => \N__44655\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44757\,
            in1 => \N__48854\,
            in2 => \_gnd_net_\,
            in3 => \N__44628\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__52399\,
            ce => 'H',
            sr => \N__51978\
        );

    \pwm_generator_inst.counter_1_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44753\,
            in1 => \N__48827\,
            in2 => \_gnd_net_\,
            in3 => \N__44625\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__52399\,
            ce => 'H',
            sr => \N__51978\
        );

    \pwm_generator_inst.counter_2_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44758\,
            in1 => \N__49382\,
            in2 => \_gnd_net_\,
            in3 => \N__44622\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__52399\,
            ce => 'H',
            sr => \N__51978\
        );

    \pwm_generator_inst.counter_3_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44754\,
            in1 => \N__49355\,
            in2 => \_gnd_net_\,
            in3 => \N__44619\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__52399\,
            ce => 'H',
            sr => \N__51978\
        );

    \pwm_generator_inst.counter_4_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44759\,
            in1 => \N__49328\,
            in2 => \_gnd_net_\,
            in3 => \N__44616\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__52399\,
            ce => 'H',
            sr => \N__51978\
        );

    \pwm_generator_inst.counter_5_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44755\,
            in1 => \N__49301\,
            in2 => \_gnd_net_\,
            in3 => \N__44613\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__52399\,
            ce => 'H',
            sr => \N__51978\
        );

    \pwm_generator_inst.counter_6_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44760\,
            in1 => \N__49271\,
            in2 => \_gnd_net_\,
            in3 => \N__44610\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__52399\,
            ce => 'H',
            sr => \N__51978\
        );

    \pwm_generator_inst.counter_7_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44756\,
            in1 => \N__49247\,
            in2 => \_gnd_net_\,
            in3 => \N__44607\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__52399\,
            ce => 'H',
            sr => \N__51978\
        );

    \pwm_generator_inst.counter_8_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44752\,
            in1 => \N__49221\,
            in2 => \_gnd_net_\,
            in3 => \N__44778\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_16_24_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__52394\,
            ce => 'H',
            sr => \N__51987\
        );

    \pwm_generator_inst.counter_9_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__49197\,
            in1 => \N__44751\,
            in2 => \_gnd_net_\,
            in3 => \N__44775\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52394\,
            ce => 'H',
            sr => \N__51987\
        );

    \pwm_generator_inst.counter_RNITBL3_9_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__49219\,
            in1 => \N__49195\,
            in2 => \_gnd_net_\,
            in3 => \N__49302\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIRPD2_0_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48855\,
            in2 => \_gnd_net_\,
            in3 => \N__48828\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_2_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__49329\,
            in1 => \N__49356\,
            in2 => \N__44772\,
            in3 => \N__49383\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_6_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__44769\,
            in1 => \N__49248\,
            in2 => \N__44763\,
            in3 => \N__49275\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100001110100"
        )
    port map (
            in0 => \N__51148\,
            in1 => \N__51369\,
            in2 => \N__44718\,
            in3 => \N__51129\,
            lcout => \pwm_generator_inst.un19_threshold_0_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__51426\,
            in1 => \N__51393\,
            in2 => \N__51379\,
            in3 => \N__51450\,
            lcout => \pwm_generator_inst.un19_threshold_0_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__51261\,
            in1 => \N__51234\,
            in2 => \N__44841\,
            in3 => \N__51367\,
            lcout => \pwm_generator_inst.un19_threshold_0_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49640\,
            in2 => \_gnd_net_\,
            in3 => \N__51191\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_16_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51221\,
            in2 => \_gnd_net_\,
            in3 => \N__45026\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_13\,
            ltout => \pwm_generator_inst.un15_threshold_1_axb_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_16_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__51368\,
            in1 => \N__51204\,
            in2 => \N__45030\,
            in3 => \N__45027\,
            lcout => \pwm_generator_inst.un19_threshold_0_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_16_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__49610\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51496\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_16_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__45012\,
            in1 => \N__45441\,
            in2 => \N__44979\,
            in3 => \N__44871\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_16_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44852\,
            in2 => \_gnd_net_\,
            in3 => \N__51080\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_17\,
            ltout => \pwm_generator_inst.un15_threshold_1_axb_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_16_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__44853\,
            in1 => \N__51370\,
            in2 => \N__44844\,
            in3 => \N__51066\,
            lcout => \pwm_generator_inst.un19_threshold_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_16_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__51115\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49664\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_16_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44834\,
            in2 => \_gnd_net_\,
            in3 => \N__51253\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_axb_4_LC_16_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44823\,
            in2 => \N__44802\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_16_28_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_16_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45357\,
            in2 => \N__45336\,
            in3 => \N__45306\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_16_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45303\,
            in2 => \N__45282\,
            in3 => \N__45255\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_16_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45252\,
            in2 => \N__45234\,
            in3 => \N__45207\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_16_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45204\,
            in2 => \N__45189\,
            in3 => \N__45168\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_16_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45165\,
            in2 => \N__45150\,
            in3 => \N__45126\,
            lcout => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_16_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45123\,
            in2 => \N__45102\,
            in3 => \N__45081\,
            lcout => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_16_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45078\,
            in2 => \N__45057\,
            in3 => \N__45033\,
            lcout => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_16_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45681\,
            in2 => \N__45660\,
            in3 => \N__45636\,
            lcout => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \bfn_16_29_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_16_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45633\,
            in2 => \N__45612\,
            in3 => \N__45585\,
            lcout => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_16_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45582\,
            in2 => \N__45438\,
            in3 => \N__45555\,
            lcout => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_16_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45426\,
            in2 => \N__45552\,
            in3 => \N__45525\,
            lcout => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_16_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45522\,
            in2 => \N__45439\,
            in3 => \N__45501\,
            lcout => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_16_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45430\,
            in2 => \N__45498\,
            in3 => \N__45474\,
            lcout => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_16_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45471\,
            in2 => \N__45440\,
            in3 => \N__45444\,
            lcout => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_16_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45434\,
            in2 => \N__45378\,
            in3 => \N__45816\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_16_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45813\,
            in1 => \N__45807\,
            in2 => \_gnd_net_\,
            in3 => \N__45798\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_red_c_g_THRU_LUT4_0_LC_16_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__52086\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_red_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_23_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46922\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52489\,
            ce => \N__50156\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45774\,
            in2 => \N__47153\,
            in3 => \N__47635\,
            lcout => \phase_controller_inst1.stoper_hc.measured_delay_hc_i_31\,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47103\,
            in1 => \N__47102\,
            in2 => \N__46757\,
            in3 => \N__45750\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_1,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47082\,
            in1 => \N__47081\,
            in2 => \N__46761\,
            in3 => \N__45726\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_2,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47058\,
            in1 => \N__47057\,
            in2 => \N__46758\,
            in3 => \N__45705\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_3,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47034\,
            in1 => \N__47033\,
            in2 => \N__46762\,
            in3 => \N__45684\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_4,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47001\,
            in1 => \N__47000\,
            in2 => \N__46759\,
            in3 => \N__45942\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_5,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__46968\,
            in1 => \N__46967\,
            in2 => \N__46763\,
            in3 => \N__45921\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_6,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47367\,
            in1 => \N__47363\,
            in2 => \N__46760\,
            in3 => \N__45903\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_7,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47334\,
            in1 => \N__47333\,
            in2 => \N__46852\,
            in3 => \N__45885\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_8,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47313\,
            in1 => \N__47312\,
            in2 => \N__46771\,
            in3 => \N__45870\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_9,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47292\,
            in1 => \N__47291\,
            in2 => \N__46853\,
            in3 => \N__45855\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_10,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47262\,
            in1 => \N__47261\,
            in2 => \N__46768\,
            in3 => \N__45837\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_11,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47235\,
            in1 => \N__47234\,
            in2 => \N__46850\,
            in3 => \N__45819\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_12,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47211\,
            in1 => \N__47210\,
            in2 => \N__46769\,
            in3 => \N__46041\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_13,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47181\,
            in1 => \N__47180\,
            in2 => \N__46851\,
            in3 => \N__46026\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_14,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47574\,
            in1 => \N__47573\,
            in2 => \N__46770\,
            in3 => \N__46011\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_15,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47541\,
            in1 => \N__47540\,
            in2 => \N__46882\,
            in3 => \N__46008\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_16,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47511\,
            in1 => \N__47510\,
            in2 => \N__46764\,
            in3 => \N__46005\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_17,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47484\,
            in1 => \N__47483\,
            in2 => \N__46883\,
            in3 => \N__46002\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_18,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47457\,
            in1 => \N__47456\,
            in2 => \N__46765\,
            in3 => \N__45999\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_19,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47436\,
            in1 => \N__47435\,
            in2 => \N__46884\,
            in3 => \N__45978\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_20,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47412\,
            in1 => \N__47411\,
            in2 => \N__46766\,
            in3 => \N__45960\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_21,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47388\,
            in1 => \N__47387\,
            in2 => \N__46885\,
            in3 => \N__46926\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_22,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47796\,
            in1 => \N__47795\,
            in2 => \N__46767\,
            in3 => \N__46899\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_23,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47775\,
            in1 => \N__47774\,
            in2 => \N__46886\,
            in3 => \N__46896\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_24,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47745\,
            in1 => \N__47744\,
            in2 => \N__46848\,
            in3 => \N__46893\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_25,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47727\,
            in1 => \N__47726\,
            in2 => \N__46887\,
            in3 => \N__46890\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_26,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47700\,
            in1 => \N__47699\,
            in2 => \N__46849\,
            in3 => \N__46101\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_27,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46098\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47625\,
            in2 => \N__46083\,
            in3 => \N__46094\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46059\,
            in2 => \_gnd_net_\,
            in3 => \N__46074\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47163\,
            in2 => \_gnd_net_\,
            in3 => \N__47115\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47112\,
            in2 => \_gnd_net_\,
            in3 => \N__47085\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50025\,
            in2 => \_gnd_net_\,
            in3 => \N__47067\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47064\,
            in2 => \_gnd_net_\,
            in3 => \N__47043\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47040\,
            in2 => \_gnd_net_\,
            in3 => \N__47016\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47013\,
            in2 => \_gnd_net_\,
            in3 => \N__46983\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46980\,
            in2 => \_gnd_net_\,
            in3 => \N__46953\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46950\,
            in2 => \_gnd_net_\,
            in3 => \N__47346\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47343\,
            in2 => \_gnd_net_\,
            in3 => \N__47316\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50031\,
            in2 => \_gnd_net_\,
            in3 => \N__47295\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50436\,
            in2 => \_gnd_net_\,
            in3 => \N__47271\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47268\,
            in2 => \_gnd_net_\,
            in3 => \N__47244\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47241\,
            in2 => \_gnd_net_\,
            in3 => \N__47220\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47217\,
            in2 => \_gnd_net_\,
            in3 => \N__47190\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47187\,
            in2 => \_gnd_net_\,
            in3 => \N__47166\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9\,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47583\,
            in2 => \_gnd_net_\,
            in3 => \N__47556\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47553\,
            in2 => \_gnd_net_\,
            in3 => \N__47523\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47520\,
            in2 => \_gnd_net_\,
            in3 => \N__47493\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47490\,
            in2 => \_gnd_net_\,
            in3 => \N__47469\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47466\,
            in2 => \_gnd_net_\,
            in3 => \N__47439\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50457\,
            in2 => \_gnd_net_\,
            in3 => \N__47421\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47418\,
            in2 => \_gnd_net_\,
            in3 => \N__47397\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47394\,
            in2 => \_gnd_net_\,
            in3 => \N__47370\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47805\,
            in2 => \_gnd_net_\,
            in3 => \N__47778\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50376\,
            in2 => \_gnd_net_\,
            in3 => \N__47760\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47757\,
            in2 => \_gnd_net_\,
            in3 => \N__47730\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50721\,
            in2 => \_gnd_net_\,
            in3 => \N__47709\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47706\,
            in2 => \_gnd_net_\,
            in3 => \N__47685\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__47682\,
            in1 => \N__47617\,
            in2 => \_gnd_net_\,
            in3 => \N__47670\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47618\,
            in1 => \N__48327\,
            in2 => \_gnd_net_\,
            in3 => \N__50835\,
            lcout => \elapsed_time_ns_1_RNI04EN9_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48299\,
            in2 => \N__50673\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__52440\,
            ce => \N__50582\,
            sr => \N__51946\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48278\,
            in2 => \N__50628\,
            in3 => \N__47586\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__52440\,
            ce => \N__50582\,
            sr => \N__51946\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48300\,
            in2 => \N__48258\,
            in3 => \N__47880\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__52440\,
            ce => \N__50582\,
            sr => \N__51946\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48279\,
            in2 => \N__48231\,
            in3 => \N__47877\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__52440\,
            ce => \N__50582\,
            sr => \N__51946\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48257\,
            in2 => \N__48197\,
            in3 => \N__47874\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__52440\,
            ce => \N__50582\,
            sr => \N__51946\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48230\,
            in2 => \N__48578\,
            in3 => \N__47871\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__52440\,
            ce => \N__50582\,
            sr => \N__51946\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48542\,
            in2 => \N__48198\,
            in3 => \N__47850\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__52440\,
            ce => \N__50582\,
            sr => \N__51946\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48512\,
            in2 => \N__48579\,
            in3 => \N__47829\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__52440\,
            ce => \N__50582\,
            sr => \N__51946\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48485\,
            in2 => \N__48549\,
            in3 => \N__47811\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__52435\,
            ce => \N__50574\,
            sr => \N__51952\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48461\,
            in2 => \N__48516\,
            in3 => \N__47808\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__52435\,
            ce => \N__50574\,
            sr => \N__51952\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48486\,
            in2 => \N__48437\,
            in3 => \N__48042\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__52435\,
            ce => \N__50574\,
            sr => \N__51952\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48462\,
            in2 => \N__48407\,
            in3 => \N__48021\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__52435\,
            ce => \N__50574\,
            sr => \N__51952\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48377\,
            in2 => \N__48438\,
            in3 => \N__48003\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__52435\,
            ce => \N__50574\,
            sr => \N__51952\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48353\,
            in2 => \N__48408\,
            in3 => \N__47982\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__52435\,
            ce => \N__50574\,
            sr => \N__51952\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48378\,
            in2 => \N__48797\,
            in3 => \N__47964\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__52435\,
            ce => \N__50574\,
            sr => \N__51952\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48354\,
            in2 => \N__48765\,
            in3 => \N__47940\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__52435\,
            ce => \N__50574\,
            sr => \N__51952\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48728\,
            in2 => \N__48798\,
            in3 => \N__47919\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__52430\,
            ce => \N__50573\,
            sr => \N__51955\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48764\,
            in2 => \N__48701\,
            in3 => \N__47898\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__52430\,
            ce => \N__50573\,
            sr => \N__51955\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48674\,
            in2 => \N__48732\,
            in3 => \N__47883\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__52430\,
            ce => \N__50573\,
            sr => \N__51955\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48650\,
            in2 => \N__48702\,
            in3 => \N__48150\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__52430\,
            ce => \N__50573\,
            sr => \N__51955\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48675\,
            in2 => \N__48626\,
            in3 => \N__48147\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__52430\,
            ce => \N__50573\,
            sr => \N__51955\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48599\,
            in2 => \N__48654\,
            in3 => \N__48126\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__52430\,
            ce => \N__50573\,
            sr => \N__51955\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49166\,
            in2 => \N__48627\,
            in3 => \N__48108\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__52430\,
            ce => \N__50573\,
            sr => \N__51955\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48600\,
            in2 => \N__49136\,
            in3 => \N__48096\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__52430\,
            ce => \N__50573\,
            sr => \N__51955\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49103\,
            in2 => \N__49173\,
            in3 => \N__48093\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__52424\,
            ce => \N__50575\,
            sr => \N__51959\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49082\,
            in2 => \N__49140\,
            in3 => \N__48069\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__52424\,
            ce => \N__50575\,
            sr => \N__51959\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49104\,
            in2 => \N__49062\,
            in3 => \N__48066\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__52424\,
            ce => \N__50575\,
            sr => \N__51959\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49083\,
            in2 => \N__48921\,
            in3 => \N__48333\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__52424\,
            ce => \N__50575\,
            sr => \N__51959\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48330\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52424\,
            ce => \N__50575\,
            sr => \N__51959\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49034\,
            in1 => \N__50662\,
            in2 => \_gnd_net_\,
            in3 => \N__48306\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__52419\,
            ce => \N__48888\,
            sr => \N__51965\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49030\,
            in1 => \N__50617\,
            in2 => \_gnd_net_\,
            in3 => \N__48303\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__52419\,
            ce => \N__48888\,
            sr => \N__51965\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49035\,
            in1 => \N__48298\,
            in2 => \_gnd_net_\,
            in3 => \N__48282\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__52419\,
            ce => \N__48888\,
            sr => \N__51965\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49031\,
            in1 => \N__48277\,
            in2 => \_gnd_net_\,
            in3 => \N__48261\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__52419\,
            ce => \N__48888\,
            sr => \N__51965\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49036\,
            in1 => \N__48253\,
            in2 => \_gnd_net_\,
            in3 => \N__48234\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__52419\,
            ce => \N__48888\,
            sr => \N__51965\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49032\,
            in1 => \N__48220\,
            in2 => \_gnd_net_\,
            in3 => \N__48201\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__52419\,
            ce => \N__48888\,
            sr => \N__51965\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49037\,
            in1 => \N__48185\,
            in2 => \_gnd_net_\,
            in3 => \N__48171\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__52419\,
            ce => \N__48888\,
            sr => \N__51965\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49033\,
            in1 => \N__48566\,
            in2 => \_gnd_net_\,
            in3 => \N__48552\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__52419\,
            ce => \N__48888\,
            sr => \N__51965\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49019\,
            in1 => \N__48541\,
            in2 => \_gnd_net_\,
            in3 => \N__48519\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__52414\,
            ce => \N__48898\,
            sr => \N__51969\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49041\,
            in1 => \N__48505\,
            in2 => \_gnd_net_\,
            in3 => \N__48489\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__52414\,
            ce => \N__48898\,
            sr => \N__51969\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49016\,
            in1 => \N__48479\,
            in2 => \_gnd_net_\,
            in3 => \N__48465\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__52414\,
            ce => \N__48898\,
            sr => \N__51969\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49038\,
            in1 => \N__48455\,
            in2 => \_gnd_net_\,
            in3 => \N__48441\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__52414\,
            ce => \N__48898\,
            sr => \N__51969\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49017\,
            in1 => \N__48425\,
            in2 => \_gnd_net_\,
            in3 => \N__48411\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__52414\,
            ce => \N__48898\,
            sr => \N__51969\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49039\,
            in1 => \N__48395\,
            in2 => \_gnd_net_\,
            in3 => \N__48381\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__52414\,
            ce => \N__48898\,
            sr => \N__51969\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49018\,
            in1 => \N__48371\,
            in2 => \_gnd_net_\,
            in3 => \N__48357\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__52414\,
            ce => \N__48898\,
            sr => \N__51969\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49040\,
            in1 => \N__48347\,
            in2 => \_gnd_net_\,
            in3 => \N__48801\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__52414\,
            ce => \N__48898\,
            sr => \N__51969\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49012\,
            in1 => \N__48784\,
            in2 => \_gnd_net_\,
            in3 => \N__48768\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__52408\,
            ce => \N__48903\,
            sr => \N__51974\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49026\,
            in1 => \N__48754\,
            in2 => \_gnd_net_\,
            in3 => \N__48735\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__52408\,
            ce => \N__48903\,
            sr => \N__51974\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49013\,
            in1 => \N__48721\,
            in2 => \_gnd_net_\,
            in3 => \N__48705\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__52408\,
            ce => \N__48903\,
            sr => \N__51974\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49027\,
            in1 => \N__48694\,
            in2 => \_gnd_net_\,
            in3 => \N__48678\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__52408\,
            ce => \N__48903\,
            sr => \N__51974\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49014\,
            in1 => \N__48673\,
            in2 => \_gnd_net_\,
            in3 => \N__48657\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__52408\,
            ce => \N__48903\,
            sr => \N__51974\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49028\,
            in1 => \N__48649\,
            in2 => \_gnd_net_\,
            in3 => \N__48630\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__52408\,
            ce => \N__48903\,
            sr => \N__51974\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49015\,
            in1 => \N__48619\,
            in2 => \_gnd_net_\,
            in3 => \N__48603\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__52408\,
            ce => \N__48903\,
            sr => \N__51974\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49029\,
            in1 => \N__48598\,
            in2 => \_gnd_net_\,
            in3 => \N__48582\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__52408\,
            ce => \N__48903\,
            sr => \N__51974\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49020\,
            in1 => \N__49165\,
            in2 => \_gnd_net_\,
            in3 => \N__49143\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_23_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__52403\,
            ce => \N__48902\,
            sr => \N__51975\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49024\,
            in1 => \N__49129\,
            in2 => \_gnd_net_\,
            in3 => \N__49107\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__52403\,
            ce => \N__48902\,
            sr => \N__51975\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49021\,
            in1 => \N__49102\,
            in2 => \_gnd_net_\,
            in3 => \N__49086\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__52403\,
            ce => \N__48902\,
            sr => \N__51975\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49025\,
            in1 => \N__49081\,
            in2 => \_gnd_net_\,
            in3 => \N__49065\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__52403\,
            ce => \N__48902\,
            sr => \N__51975\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49022\,
            in1 => \N__49058\,
            in2 => \_gnd_net_\,
            in3 => \N__49044\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__52403\,
            ce => \N__48902\,
            sr => \N__51975\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__48917\,
            in1 => \N__49023\,
            in2 => \_gnd_net_\,
            in3 => \N__48924\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52403\,
            ce => \N__48902\,
            sr => \N__51975\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__48853\,
            in1 => \N__48834\,
            in2 => \N__49524\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_17_24_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48807\,
            in2 => \N__49509\,
            in3 => \N__48826\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49362\,
            in2 => \N__49482\,
            in3 => \N__49378\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__49351\,
            in1 => \N__49335\,
            in2 => \N__49458\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__49324\,
            in1 => \N__49308\,
            in2 => \N__49440\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49281\,
            in2 => \N__49419\,
            in3 => \N__49297\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49254\,
            in2 => \N__49401\,
            in3 => \N__49270\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__49243\,
            in1 => \N__49227\,
            in2 => \N__49731\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__49220\,
            in1 => \N__49203\,
            in2 => \N__49713\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_17_25_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49179\,
            in2 => \N__49683\,
            in3 => \N__49196\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49557\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52395\,
            ce => 'H',
            sr => \N__51988\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_17_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49530\,
            in2 => \N__51381\,
            in3 => \N__51380\,
            lcout => \pwm_generator_inst.un14_counter_0\,
            ltout => OPEN,
            carryin => \bfn_17_26_0_\,
            carryout => \pwm_generator_inst.un19_threshold_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_0_cry_0_c_RNI2C682_LC_17_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51273\,
            in2 => \_gnd_net_\,
            in3 => \N__49494\,
            lcout => \pwm_generator_inst.un14_counter_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_0_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_0_cry_1_c_RNI93892_LC_17_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__49491\,
            in3 => \N__49467\,
            lcout => \pwm_generator_inst.un14_counter_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_0_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_0_cry_2_c_RNIC9B92_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49464\,
            in2 => \_gnd_net_\,
            in3 => \N__49443\,
            lcout => \pwm_generator_inst.un14_counter_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_0_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_0_cry_3_c_RNIFFE92_LC_17_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49623\,
            in2 => \_gnd_net_\,
            in3 => \N__49428\,
            lcout => \pwm_generator_inst.un14_counter_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_0_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_0_cry_4_c_RNI0V9N2_LC_17_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49425\,
            in2 => \_gnd_net_\,
            in3 => \N__49404\,
            lcout => \pwm_generator_inst.un14_counter_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_0_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_0_cry_5_c_RNIVCMU2_LC_17_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49653\,
            in2 => \_gnd_net_\,
            in3 => \N__49386\,
            lcout => \pwm_generator_inst.un14_counter_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_0_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_0_cry_6_c_RNI3LQU2_LC_17_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49737\,
            in2 => \_gnd_net_\,
            in3 => \N__49716\,
            lcout => \pwm_generator_inst.un14_counter_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_0_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_0_cry_7_c_RNI7TUU2_LC_17_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49599\,
            in2 => \_gnd_net_\,
            in3 => \N__49701\,
            lcout => \pwm_generator_inst.un14_counter_8\,
            ltout => OPEN,
            carryin => \bfn_17_27_0_\,
            carryout => \pwm_generator_inst.un19_threshold_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIB53V2_LC_17_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__51459\,
            in1 => \N__49698\,
            in2 => \N__51378\,
            in3 => \N__49686\,
            lcout => \pwm_generator_inst.un14_counter_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_17_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011110000100"
        )
    port map (
            in0 => \N__51093\,
            in1 => \N__51359\,
            in2 => \N__51117\,
            in3 => \N__49671\,
            lcout => \pwm_generator_inst.un19_threshold_0_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_17_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__51171\,
            in1 => \N__51190\,
            in2 => \N__49647\,
            in3 => \N__51358\,
            lcout => \pwm_generator_inst.un19_threshold_0_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_17_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__51360\,
            in1 => \N__49617\,
            in2 => \N__51498\,
            in3 => \N__51474\,
            lcout => \pwm_generator_inst.un19_threshold_0_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_16_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49593\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52490\,
            ce => \N__50141\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_18_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49577\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52490\,
            ce => \N__50141\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_19_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50019\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52490\,
            ce => \N__50141\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__49992\,
            in1 => \N__49982\,
            in2 => \N__49964\,
            in3 => \N__49905\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__49991\,
            in1 => \N__49983\,
            in2 => \N__49965\,
            in3 => \N__49904\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_17_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49916\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52484\,
            ce => \N__50157\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__49881\,
            in1 => \N__49872\,
            in2 => \N__49850\,
            in3 => \N__49827\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__49880\,
            in1 => \N__49871\,
            in2 => \N__49851\,
            in3 => \N__49826\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__50193\,
            in1 => \N__49791\,
            in2 => \N__50172\,
            in3 => \N__49773\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__50192\,
            in1 => \N__49790\,
            in2 => \N__50171\,
            in3 => \N__49772\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__50214\,
            in1 => \N__50307\,
            in2 => \N__50288\,
            in3 => \N__50235\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__50213\,
            in1 => \N__50306\,
            in2 => \N__50289\,
            in3 => \N__50234\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_27_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50247\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52481\,
            ce => \N__50140\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_26_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50226\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52477\,
            ce => \N__50148\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_24_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50205\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52477\,
            ce => \N__50148\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_25_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50184\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52477\,
            ce => \N__50148\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50040\,
            in1 => \N__50061\,
            in2 => \_gnd_net_\,
            in3 => \N__50875\,
            lcout => \elapsed_time_ns_1_RNIV0CN9_0_12\,
            ltout => \elapsed_time_ns_1_RNIV0CN9_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50034\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__50447\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50466\,
            in1 => \N__50484\,
            in2 => \_gnd_net_\,
            in3 => \N__50876\,
            lcout => \elapsed_time_ns_1_RNI14DN9_0_23\,
            ltout => \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50460\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50358\,
            in1 => \N__50448\,
            in2 => \_gnd_net_\,
            in3 => \N__50874\,
            lcout => \elapsed_time_ns_1_RNIH33T9_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50414\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50877\,
            in1 => \N__50415\,
            in2 => \_gnd_net_\,
            in3 => \N__50430\,
            lcout => \elapsed_time_ns_1_RNI02CN9_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50385\,
            in1 => \N__50403\,
            in2 => \_gnd_net_\,
            in3 => \N__50878\,
            lcout => \elapsed_time_ns_1_RNI58DN9_0_27\,
            ltout => \elapsed_time_ns_1_RNI58DN9_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50379\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50369\,
            in2 => \_gnd_net_\,
            in3 => \N__50354\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__50336\,
            in1 => \N__50321\,
            in2 => \N__50310\,
            in3 => \N__50679\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50730\,
            in1 => \N__50898\,
            in2 => \_gnd_net_\,
            in3 => \N__50879\,
            lcout => \elapsed_time_ns_1_RNI7ADN9_0_29\,
            ltout => \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50724\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__50708\,
            in1 => \N__50594\,
            in2 => \N__50696\,
            in3 => \N__50639\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50672\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52447\,
            ce => \N__50583\,
            sr => \N__51944\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50627\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52447\,
            ce => \N__50583\,
            sr => \N__51944\
        );

    \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_20_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50526\,
            in2 => \_gnd_net_\,
            in3 => \N__50541\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_20_25_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_20_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50508\,
            in2 => \_gnd_net_\,
            in3 => \N__50520\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_20_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50490\,
            in2 => \_gnd_net_\,
            in3 => \N__50502\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_20_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51036\,
            in2 => \_gnd_net_\,
            in3 => \N__51051\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_20_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51015\,
            in2 => \_gnd_net_\,
            in3 => \N__51030\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_20_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50994\,
            in2 => \_gnd_net_\,
            in3 => \N__51009\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_20_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50973\,
            in2 => \_gnd_net_\,
            in3 => \N__50988\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_20_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50952\,
            in2 => \_gnd_net_\,
            in3 => \N__50967\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_20_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50931\,
            in2 => \_gnd_net_\,
            in3 => \N__50946\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_20_26_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_20_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50913\,
            in2 => \_gnd_net_\,
            in3 => \N__50925\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_20_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51421\,
            in2 => \_gnd_net_\,
            in3 => \N__51384\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_20_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__51374\,
            in1 => \N__51299\,
            in2 => \_gnd_net_\,
            in3 => \N__51264\,
            lcout => \pwm_generator_inst.un19_threshold_0_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_20_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51260\,
            in2 => \_gnd_net_\,
            in3 => \N__51225\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_20_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51222\,
            in2 => \_gnd_net_\,
            in3 => \N__51195\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_20_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51192\,
            in2 => \_gnd_net_\,
            in3 => \N__51159\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_20_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51156\,
            in2 => \_gnd_net_\,
            in3 => \N__51120\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_20_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51116\,
            in2 => \_gnd_net_\,
            in3 => \N__51084\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_20_27_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_20_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51081\,
            in2 => \_gnd_net_\,
            in3 => \N__51054\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_20_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51497\,
            in2 => \_gnd_net_\,
            in3 => \N__51465\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_20_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51462\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_21_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__52726\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52825\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_21_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__51425\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51449\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_22_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52774\,
            in2 => \_gnd_net_\,
            in3 => \N__52727\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52862\,
            in1 => \N__51405\,
            in2 => \N__52826\,
            in3 => \N__52532\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__52531\,
            in1 => \N__52861\,
            in2 => \N__52781\,
            in3 => \N__51399\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52929\,
            in2 => \_gnd_net_\,
            in3 => \N__51562\,
            lcout => \current_shift_inst.PI_CTRL.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__52625\,
            in1 => \N__51676\,
            in2 => \N__52939\,
            in3 => \N__52561\,
            lcout => \current_shift_inst.PI_CTRL.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_23_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__51693\,
            in1 => \N__52626\,
            in2 => \N__52895\,
            in3 => \N__52672\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => \current_shift_inst.PI_CTRL.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_23_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__51563\,
            in1 => \N__51684\,
            in2 => \N__51687\,
            in3 => \N__51527\,
            lcout => \current_shift_inst.PI_CTRL.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__51677\,
            in1 => \N__52560\,
            in2 => \_gnd_net_\,
            in3 => \N__52624\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__52627\,
            in1 => \N__51678\,
            in2 => \N__52940\,
            in3 => \N__52562\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_24_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51666\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52454\,
            ce => 'H',
            sr => \N__51979\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_24_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__51606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51651\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52448\,
            ce => 'H',
            sr => \N__51990\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__51621\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51604\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52448\,
            ce => 'H',
            sr => \N__51990\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_24_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__51605\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51594\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52448\,
            ce => 'H',
            sr => \N__51990\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__51567\,
            in1 => \N__51528\,
            in2 => \_gnd_net_\,
            in3 => \N__51516\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52448\,
            ce => 'H',
            sr => \N__51990\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010101010101"
        )
    port map (
            in0 => \N__52947\,
            in1 => \N__52941\,
            in2 => \N__52899\,
            in3 => \N__52692\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52448\,
            ce => 'H',
            sr => \N__51990\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__52650\,
            in1 => \N__52691\,
            in2 => \N__52869\,
            in3 => \N__52587\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52441\,
            ce => 'H',
            sr => \N__51994\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110000"
        )
    port map (
            in0 => \N__52688\,
            in1 => \N__52647\,
            in2 => \N__52588\,
            in3 => \N__52827\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52441\,
            ce => 'H',
            sr => \N__51994\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_24_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__52646\,
            in1 => \N__52687\,
            in2 => \N__52782\,
            in3 => \N__52586\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52441\,
            ce => 'H',
            sr => \N__51994\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110000"
        )
    port map (
            in0 => \N__52690\,
            in1 => \N__52649\,
            in2 => \N__52590\,
            in3 => \N__52731\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52441\,
            ce => 'H',
            sr => \N__51994\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_24_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110000"
        )
    port map (
            in0 => \N__52689\,
            in1 => \N__52648\,
            in2 => \N__52589\,
            in3 => \N__52536\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52441\,
            ce => 'H',
            sr => \N__51994\
        );
end \INTERFACE\;
