-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Oct 3 2024 21:46:45

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    start_stop : in std_logic;
    s2_phy : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    error_pin : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__54407\ : std_logic;
signal \N__54406\ : std_logic;
signal \N__54405\ : std_logic;
signal \N__54396\ : std_logic;
signal \N__54395\ : std_logic;
signal \N__54394\ : std_logic;
signal \N__54387\ : std_logic;
signal \N__54386\ : std_logic;
signal \N__54385\ : std_logic;
signal \N__54378\ : std_logic;
signal \N__54377\ : std_logic;
signal \N__54376\ : std_logic;
signal \N__54369\ : std_logic;
signal \N__54368\ : std_logic;
signal \N__54367\ : std_logic;
signal \N__54360\ : std_logic;
signal \N__54359\ : std_logic;
signal \N__54358\ : std_logic;
signal \N__54351\ : std_logic;
signal \N__54350\ : std_logic;
signal \N__54349\ : std_logic;
signal \N__54342\ : std_logic;
signal \N__54341\ : std_logic;
signal \N__54340\ : std_logic;
signal \N__54333\ : std_logic;
signal \N__54332\ : std_logic;
signal \N__54331\ : std_logic;
signal \N__54324\ : std_logic;
signal \N__54323\ : std_logic;
signal \N__54322\ : std_logic;
signal \N__54315\ : std_logic;
signal \N__54314\ : std_logic;
signal \N__54313\ : std_logic;
signal \N__54306\ : std_logic;
signal \N__54305\ : std_logic;
signal \N__54304\ : std_logic;
signal \N__54297\ : std_logic;
signal \N__54296\ : std_logic;
signal \N__54295\ : std_logic;
signal \N__54278\ : std_logic;
signal \N__54275\ : std_logic;
signal \N__54274\ : std_logic;
signal \N__54269\ : std_logic;
signal \N__54266\ : std_logic;
signal \N__54263\ : std_logic;
signal \N__54262\ : std_logic;
signal \N__54261\ : std_logic;
signal \N__54260\ : std_logic;
signal \N__54259\ : std_logic;
signal \N__54252\ : std_logic;
signal \N__54249\ : std_logic;
signal \N__54248\ : std_logic;
signal \N__54247\ : std_logic;
signal \N__54246\ : std_logic;
signal \N__54243\ : std_logic;
signal \N__54240\ : std_logic;
signal \N__54237\ : std_logic;
signal \N__54232\ : std_logic;
signal \N__54229\ : std_logic;
signal \N__54222\ : std_logic;
signal \N__54217\ : std_logic;
signal \N__54214\ : std_logic;
signal \N__54211\ : std_logic;
signal \N__54208\ : std_logic;
signal \N__54205\ : std_logic;
signal \N__54202\ : std_logic;
signal \N__54199\ : std_logic;
signal \N__54194\ : std_logic;
signal \N__54191\ : std_logic;
signal \N__54190\ : std_logic;
signal \N__54187\ : std_logic;
signal \N__54184\ : std_logic;
signal \N__54179\ : std_logic;
signal \N__54178\ : std_logic;
signal \N__54177\ : std_logic;
signal \N__54170\ : std_logic;
signal \N__54167\ : std_logic;
signal \N__54166\ : std_logic;
signal \N__54165\ : std_logic;
signal \N__54164\ : std_logic;
signal \N__54161\ : std_logic;
signal \N__54158\ : std_logic;
signal \N__54155\ : std_logic;
signal \N__54152\ : std_logic;
signal \N__54147\ : std_logic;
signal \N__54144\ : std_logic;
signal \N__54141\ : std_logic;
signal \N__54138\ : std_logic;
signal \N__54133\ : std_logic;
signal \N__54130\ : std_logic;
signal \N__54127\ : std_logic;
signal \N__54124\ : std_logic;
signal \N__54121\ : std_logic;
signal \N__54116\ : std_logic;
signal \N__54115\ : std_logic;
signal \N__54114\ : std_logic;
signal \N__54111\ : std_logic;
signal \N__54108\ : std_logic;
signal \N__54105\ : std_logic;
signal \N__54098\ : std_logic;
signal \N__54095\ : std_logic;
signal \N__54092\ : std_logic;
signal \N__54091\ : std_logic;
signal \N__54090\ : std_logic;
signal \N__54089\ : std_logic;
signal \N__54088\ : std_logic;
signal \N__54087\ : std_logic;
signal \N__54086\ : std_logic;
signal \N__54085\ : std_logic;
signal \N__54080\ : std_logic;
signal \N__54073\ : std_logic;
signal \N__54068\ : std_logic;
signal \N__54067\ : std_logic;
signal \N__54064\ : std_logic;
signal \N__54063\ : std_logic;
signal \N__54056\ : std_logic;
signal \N__54053\ : std_logic;
signal \N__54050\ : std_logic;
signal \N__54047\ : std_logic;
signal \N__54042\ : std_logic;
signal \N__54037\ : std_logic;
signal \N__54034\ : std_logic;
signal \N__54031\ : std_logic;
signal \N__54028\ : std_logic;
signal \N__54025\ : std_logic;
signal \N__54022\ : std_logic;
signal \N__54019\ : std_logic;
signal \N__54014\ : std_logic;
signal \N__54011\ : std_logic;
signal \N__54010\ : std_logic;
signal \N__54007\ : std_logic;
signal \N__54004\ : std_logic;
signal \N__53999\ : std_logic;
signal \N__53996\ : std_logic;
signal \N__53995\ : std_logic;
signal \N__53994\ : std_logic;
signal \N__53993\ : std_logic;
signal \N__53992\ : std_logic;
signal \N__53989\ : std_logic;
signal \N__53986\ : std_logic;
signal \N__53983\ : std_logic;
signal \N__53982\ : std_logic;
signal \N__53979\ : std_logic;
signal \N__53976\ : std_logic;
signal \N__53973\ : std_logic;
signal \N__53966\ : std_logic;
signal \N__53965\ : std_logic;
signal \N__53960\ : std_logic;
signal \N__53957\ : std_logic;
signal \N__53954\ : std_logic;
signal \N__53951\ : std_logic;
signal \N__53948\ : std_logic;
signal \N__53943\ : std_logic;
signal \N__53940\ : std_logic;
signal \N__53937\ : std_logic;
signal \N__53934\ : std_logic;
signal \N__53931\ : std_logic;
signal \N__53928\ : std_logic;
signal \N__53925\ : std_logic;
signal \N__53922\ : std_logic;
signal \N__53915\ : std_logic;
signal \N__53912\ : std_logic;
signal \N__53911\ : std_logic;
signal \N__53908\ : std_logic;
signal \N__53905\ : std_logic;
signal \N__53900\ : std_logic;
signal \N__53897\ : std_logic;
signal \N__53894\ : std_logic;
signal \N__53891\ : std_logic;
signal \N__53890\ : std_logic;
signal \N__53887\ : std_logic;
signal \N__53884\ : std_logic;
signal \N__53881\ : std_logic;
signal \N__53878\ : std_logic;
signal \N__53875\ : std_logic;
signal \N__53872\ : std_logic;
signal \N__53869\ : std_logic;
signal \N__53864\ : std_logic;
signal \N__53861\ : std_logic;
signal \N__53858\ : std_logic;
signal \N__53855\ : std_logic;
signal \N__53854\ : std_logic;
signal \N__53853\ : std_logic;
signal \N__53852\ : std_logic;
signal \N__53851\ : std_logic;
signal \N__53850\ : std_logic;
signal \N__53849\ : std_logic;
signal \N__53848\ : std_logic;
signal \N__53847\ : std_logic;
signal \N__53846\ : std_logic;
signal \N__53845\ : std_logic;
signal \N__53844\ : std_logic;
signal \N__53843\ : std_logic;
signal \N__53842\ : std_logic;
signal \N__53841\ : std_logic;
signal \N__53840\ : std_logic;
signal \N__53839\ : std_logic;
signal \N__53838\ : std_logic;
signal \N__53837\ : std_logic;
signal \N__53836\ : std_logic;
signal \N__53835\ : std_logic;
signal \N__53834\ : std_logic;
signal \N__53833\ : std_logic;
signal \N__53832\ : std_logic;
signal \N__53831\ : std_logic;
signal \N__53830\ : std_logic;
signal \N__53829\ : std_logic;
signal \N__53828\ : std_logic;
signal \N__53827\ : std_logic;
signal \N__53826\ : std_logic;
signal \N__53825\ : std_logic;
signal \N__53824\ : std_logic;
signal \N__53823\ : std_logic;
signal \N__53822\ : std_logic;
signal \N__53821\ : std_logic;
signal \N__53820\ : std_logic;
signal \N__53819\ : std_logic;
signal \N__53818\ : std_logic;
signal \N__53817\ : std_logic;
signal \N__53816\ : std_logic;
signal \N__53815\ : std_logic;
signal \N__53814\ : std_logic;
signal \N__53813\ : std_logic;
signal \N__53812\ : std_logic;
signal \N__53811\ : std_logic;
signal \N__53810\ : std_logic;
signal \N__53809\ : std_logic;
signal \N__53808\ : std_logic;
signal \N__53807\ : std_logic;
signal \N__53806\ : std_logic;
signal \N__53805\ : std_logic;
signal \N__53804\ : std_logic;
signal \N__53803\ : std_logic;
signal \N__53802\ : std_logic;
signal \N__53801\ : std_logic;
signal \N__53800\ : std_logic;
signal \N__53799\ : std_logic;
signal \N__53798\ : std_logic;
signal \N__53797\ : std_logic;
signal \N__53796\ : std_logic;
signal \N__53795\ : std_logic;
signal \N__53794\ : std_logic;
signal \N__53793\ : std_logic;
signal \N__53792\ : std_logic;
signal \N__53791\ : std_logic;
signal \N__53790\ : std_logic;
signal \N__53789\ : std_logic;
signal \N__53788\ : std_logic;
signal \N__53787\ : std_logic;
signal \N__53786\ : std_logic;
signal \N__53785\ : std_logic;
signal \N__53784\ : std_logic;
signal \N__53783\ : std_logic;
signal \N__53782\ : std_logic;
signal \N__53781\ : std_logic;
signal \N__53780\ : std_logic;
signal \N__53779\ : std_logic;
signal \N__53778\ : std_logic;
signal \N__53777\ : std_logic;
signal \N__53776\ : std_logic;
signal \N__53775\ : std_logic;
signal \N__53774\ : std_logic;
signal \N__53773\ : std_logic;
signal \N__53772\ : std_logic;
signal \N__53771\ : std_logic;
signal \N__53770\ : std_logic;
signal \N__53769\ : std_logic;
signal \N__53768\ : std_logic;
signal \N__53767\ : std_logic;
signal \N__53766\ : std_logic;
signal \N__53765\ : std_logic;
signal \N__53764\ : std_logic;
signal \N__53763\ : std_logic;
signal \N__53762\ : std_logic;
signal \N__53761\ : std_logic;
signal \N__53760\ : std_logic;
signal \N__53759\ : std_logic;
signal \N__53758\ : std_logic;
signal \N__53757\ : std_logic;
signal \N__53756\ : std_logic;
signal \N__53755\ : std_logic;
signal \N__53754\ : std_logic;
signal \N__53753\ : std_logic;
signal \N__53752\ : std_logic;
signal \N__53751\ : std_logic;
signal \N__53750\ : std_logic;
signal \N__53749\ : std_logic;
signal \N__53748\ : std_logic;
signal \N__53747\ : std_logic;
signal \N__53746\ : std_logic;
signal \N__53745\ : std_logic;
signal \N__53744\ : std_logic;
signal \N__53743\ : std_logic;
signal \N__53742\ : std_logic;
signal \N__53741\ : std_logic;
signal \N__53740\ : std_logic;
signal \N__53739\ : std_logic;
signal \N__53738\ : std_logic;
signal \N__53737\ : std_logic;
signal \N__53736\ : std_logic;
signal \N__53735\ : std_logic;
signal \N__53734\ : std_logic;
signal \N__53733\ : std_logic;
signal \N__53732\ : std_logic;
signal \N__53731\ : std_logic;
signal \N__53730\ : std_logic;
signal \N__53729\ : std_logic;
signal \N__53728\ : std_logic;
signal \N__53727\ : std_logic;
signal \N__53468\ : std_logic;
signal \N__53465\ : std_logic;
signal \N__53464\ : std_logic;
signal \N__53463\ : std_logic;
signal \N__53462\ : std_logic;
signal \N__53461\ : std_logic;
signal \N__53460\ : std_logic;
signal \N__53459\ : std_logic;
signal \N__53458\ : std_logic;
signal \N__53455\ : std_logic;
signal \N__53452\ : std_logic;
signal \N__53449\ : std_logic;
signal \N__53446\ : std_logic;
signal \N__53443\ : std_logic;
signal \N__53440\ : std_logic;
signal \N__53437\ : std_logic;
signal \N__53434\ : std_logic;
signal \N__53431\ : std_logic;
signal \N__53428\ : std_logic;
signal \N__53425\ : std_logic;
signal \N__53424\ : std_logic;
signal \N__53423\ : std_logic;
signal \N__53422\ : std_logic;
signal \N__53419\ : std_logic;
signal \N__53418\ : std_logic;
signal \N__53417\ : std_logic;
signal \N__53416\ : std_logic;
signal \N__53415\ : std_logic;
signal \N__53414\ : std_logic;
signal \N__53413\ : std_logic;
signal \N__53412\ : std_logic;
signal \N__53411\ : std_logic;
signal \N__53410\ : std_logic;
signal \N__53409\ : std_logic;
signal \N__53408\ : std_logic;
signal \N__53407\ : std_logic;
signal \N__53406\ : std_logic;
signal \N__53405\ : std_logic;
signal \N__53404\ : std_logic;
signal \N__53403\ : std_logic;
signal \N__53402\ : std_logic;
signal \N__53401\ : std_logic;
signal \N__53400\ : std_logic;
signal \N__53397\ : std_logic;
signal \N__53396\ : std_logic;
signal \N__53395\ : std_logic;
signal \N__53394\ : std_logic;
signal \N__53393\ : std_logic;
signal \N__53392\ : std_logic;
signal \N__53391\ : std_logic;
signal \N__53390\ : std_logic;
signal \N__53389\ : std_logic;
signal \N__53388\ : std_logic;
signal \N__53387\ : std_logic;
signal \N__53386\ : std_logic;
signal \N__53385\ : std_logic;
signal \N__53384\ : std_logic;
signal \N__53383\ : std_logic;
signal \N__53382\ : std_logic;
signal \N__53381\ : std_logic;
signal \N__53380\ : std_logic;
signal \N__53379\ : std_logic;
signal \N__53378\ : std_logic;
signal \N__53377\ : std_logic;
signal \N__53376\ : std_logic;
signal \N__53375\ : std_logic;
signal \N__53374\ : std_logic;
signal \N__53373\ : std_logic;
signal \N__53372\ : std_logic;
signal \N__53371\ : std_logic;
signal \N__53370\ : std_logic;
signal \N__53369\ : std_logic;
signal \N__53368\ : std_logic;
signal \N__53367\ : std_logic;
signal \N__53366\ : std_logic;
signal \N__53365\ : std_logic;
signal \N__53364\ : std_logic;
signal \N__53363\ : std_logic;
signal \N__53362\ : std_logic;
signal \N__53359\ : std_logic;
signal \N__53358\ : std_logic;
signal \N__53357\ : std_logic;
signal \N__53356\ : std_logic;
signal \N__53355\ : std_logic;
signal \N__53354\ : std_logic;
signal \N__53351\ : std_logic;
signal \N__53350\ : std_logic;
signal \N__53349\ : std_logic;
signal \N__53348\ : std_logic;
signal \N__53347\ : std_logic;
signal \N__53346\ : std_logic;
signal \N__53345\ : std_logic;
signal \N__53344\ : std_logic;
signal \N__53343\ : std_logic;
signal \N__53342\ : std_logic;
signal \N__53341\ : std_logic;
signal \N__53340\ : std_logic;
signal \N__53339\ : std_logic;
signal \N__53338\ : std_logic;
signal \N__53337\ : std_logic;
signal \N__53336\ : std_logic;
signal \N__53335\ : std_logic;
signal \N__53332\ : std_logic;
signal \N__53331\ : std_logic;
signal \N__53330\ : std_logic;
signal \N__53329\ : std_logic;
signal \N__53328\ : std_logic;
signal \N__53327\ : std_logic;
signal \N__53326\ : std_logic;
signal \N__53325\ : std_logic;
signal \N__53324\ : std_logic;
signal \N__53323\ : std_logic;
signal \N__53322\ : std_logic;
signal \N__53321\ : std_logic;
signal \N__53320\ : std_logic;
signal \N__53319\ : std_logic;
signal \N__53318\ : std_logic;
signal \N__53317\ : std_logic;
signal \N__53316\ : std_logic;
signal \N__53315\ : std_logic;
signal \N__53314\ : std_logic;
signal \N__53313\ : std_logic;
signal \N__53312\ : std_logic;
signal \N__53099\ : std_logic;
signal \N__53096\ : std_logic;
signal \N__53093\ : std_logic;
signal \N__53092\ : std_logic;
signal \N__53091\ : std_logic;
signal \N__53086\ : std_logic;
signal \N__53083\ : std_logic;
signal \N__53080\ : std_logic;
signal \N__53077\ : std_logic;
signal \N__53074\ : std_logic;
signal \N__53071\ : std_logic;
signal \N__53068\ : std_logic;
signal \N__53063\ : std_logic;
signal \N__53060\ : std_logic;
signal \N__53057\ : std_logic;
signal \N__53056\ : std_logic;
signal \N__53053\ : std_logic;
signal \N__53050\ : std_logic;
signal \N__53047\ : std_logic;
signal \N__53044\ : std_logic;
signal \N__53043\ : std_logic;
signal \N__53040\ : std_logic;
signal \N__53037\ : std_logic;
signal \N__53034\ : std_logic;
signal \N__53031\ : std_logic;
signal \N__53026\ : std_logic;
signal \N__53023\ : std_logic;
signal \N__53020\ : std_logic;
signal \N__53017\ : std_logic;
signal \N__53014\ : std_logic;
signal \N__53009\ : std_logic;
signal \N__53006\ : std_logic;
signal \N__53003\ : std_logic;
signal \N__53002\ : std_logic;
signal \N__52999\ : std_logic;
signal \N__52996\ : std_logic;
signal \N__52993\ : std_logic;
signal \N__52990\ : std_logic;
signal \N__52989\ : std_logic;
signal \N__52984\ : std_logic;
signal \N__52981\ : std_logic;
signal \N__52976\ : std_logic;
signal \N__52973\ : std_logic;
signal \N__52970\ : std_logic;
signal \N__52967\ : std_logic;
signal \N__52964\ : std_logic;
signal \N__52961\ : std_logic;
signal \N__52958\ : std_logic;
signal \N__52955\ : std_logic;
signal \N__52952\ : std_logic;
signal \N__52949\ : std_logic;
signal \N__52946\ : std_logic;
signal \N__52943\ : std_logic;
signal \N__52940\ : std_logic;
signal \N__52937\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52931\ : std_logic;
signal \N__52928\ : std_logic;
signal \N__52925\ : std_logic;
signal \N__52922\ : std_logic;
signal \N__52919\ : std_logic;
signal \N__52916\ : std_logic;
signal \N__52913\ : std_logic;
signal \N__52910\ : std_logic;
signal \N__52907\ : std_logic;
signal \N__52904\ : std_logic;
signal \N__52901\ : std_logic;
signal \N__52898\ : std_logic;
signal \N__52895\ : std_logic;
signal \N__52892\ : std_logic;
signal \N__52889\ : std_logic;
signal \N__52886\ : std_logic;
signal \N__52883\ : std_logic;
signal \N__52880\ : std_logic;
signal \N__52877\ : std_logic;
signal \N__52874\ : std_logic;
signal \N__52871\ : std_logic;
signal \N__52868\ : std_logic;
signal \N__52865\ : std_logic;
signal \N__52862\ : std_logic;
signal \N__52859\ : std_logic;
signal \N__52856\ : std_logic;
signal \N__52853\ : std_logic;
signal \N__52850\ : std_logic;
signal \N__52847\ : std_logic;
signal \N__52844\ : std_logic;
signal \N__52841\ : std_logic;
signal \N__52838\ : std_logic;
signal \N__52835\ : std_logic;
signal \N__52832\ : std_logic;
signal \N__52831\ : std_logic;
signal \N__52830\ : std_logic;
signal \N__52827\ : std_logic;
signal \N__52824\ : std_logic;
signal \N__52821\ : std_logic;
signal \N__52814\ : std_logic;
signal \N__52811\ : std_logic;
signal \N__52808\ : std_logic;
signal \N__52805\ : std_logic;
signal \N__52802\ : std_logic;
signal \N__52799\ : std_logic;
signal \N__52796\ : std_logic;
signal \N__52795\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52793\ : std_logic;
signal \N__52792\ : std_logic;
signal \N__52791\ : std_logic;
signal \N__52790\ : std_logic;
signal \N__52789\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52787\ : std_logic;
signal \N__52786\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52784\ : std_logic;
signal \N__52783\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52781\ : std_logic;
signal \N__52764\ : std_logic;
signal \N__52747\ : std_logic;
signal \N__52742\ : std_logic;
signal \N__52739\ : std_logic;
signal \N__52738\ : std_logic;
signal \N__52737\ : std_logic;
signal \N__52736\ : std_logic;
signal \N__52735\ : std_logic;
signal \N__52734\ : std_logic;
signal \N__52731\ : std_logic;
signal \N__52726\ : std_logic;
signal \N__52719\ : std_logic;
signal \N__52716\ : std_logic;
signal \N__52711\ : std_logic;
signal \N__52708\ : std_logic;
signal \N__52703\ : std_logic;
signal \N__52700\ : std_logic;
signal \N__52699\ : std_logic;
signal \N__52698\ : std_logic;
signal \N__52695\ : std_logic;
signal \N__52690\ : std_logic;
signal \N__52687\ : std_logic;
signal \N__52684\ : std_logic;
signal \N__52681\ : std_logic;
signal \N__52678\ : std_logic;
signal \N__52675\ : std_logic;
signal \N__52672\ : std_logic;
signal \N__52667\ : std_logic;
signal \N__52664\ : std_logic;
signal \N__52661\ : std_logic;
signal \N__52658\ : std_logic;
signal \N__52655\ : std_logic;
signal \N__52652\ : std_logic;
signal \N__52649\ : std_logic;
signal \N__52648\ : std_logic;
signal \N__52643\ : std_logic;
signal \N__52640\ : std_logic;
signal \N__52637\ : std_logic;
signal \N__52634\ : std_logic;
signal \N__52631\ : std_logic;
signal \N__52628\ : std_logic;
signal \N__52625\ : std_logic;
signal \N__52622\ : std_logic;
signal \N__52621\ : std_logic;
signal \N__52618\ : std_logic;
signal \N__52615\ : std_logic;
signal \N__52612\ : std_logic;
signal \N__52609\ : std_logic;
signal \N__52606\ : std_logic;
signal \N__52601\ : std_logic;
signal \N__52600\ : std_logic;
signal \N__52597\ : std_logic;
signal \N__52594\ : std_logic;
signal \N__52591\ : std_logic;
signal \N__52588\ : std_logic;
signal \N__52585\ : std_logic;
signal \N__52580\ : std_logic;
signal \N__52579\ : std_logic;
signal \N__52576\ : std_logic;
signal \N__52573\ : std_logic;
signal \N__52570\ : std_logic;
signal \N__52567\ : std_logic;
signal \N__52564\ : std_logic;
signal \N__52559\ : std_logic;
signal \N__52558\ : std_logic;
signal \N__52555\ : std_logic;
signal \N__52550\ : std_logic;
signal \N__52547\ : std_logic;
signal \N__52544\ : std_logic;
signal \N__52543\ : std_logic;
signal \N__52538\ : std_logic;
signal \N__52535\ : std_logic;
signal \N__52532\ : std_logic;
signal \N__52531\ : std_logic;
signal \N__52526\ : std_logic;
signal \N__52523\ : std_logic;
signal \N__52520\ : std_logic;
signal \N__52519\ : std_logic;
signal \N__52514\ : std_logic;
signal \N__52511\ : std_logic;
signal \N__52508\ : std_logic;
signal \N__52505\ : std_logic;
signal \N__52504\ : std_logic;
signal \N__52501\ : std_logic;
signal \N__52498\ : std_logic;
signal \N__52495\ : std_logic;
signal \N__52490\ : std_logic;
signal \N__52487\ : std_logic;
signal \N__52484\ : std_logic;
signal \N__52481\ : std_logic;
signal \N__52478\ : std_logic;
signal \N__52475\ : std_logic;
signal \N__52472\ : std_logic;
signal \N__52469\ : std_logic;
signal \N__52466\ : std_logic;
signal \N__52463\ : std_logic;
signal \N__52462\ : std_logic;
signal \N__52459\ : std_logic;
signal \N__52456\ : std_logic;
signal \N__52455\ : std_logic;
signal \N__52454\ : std_logic;
signal \N__52451\ : std_logic;
signal \N__52448\ : std_logic;
signal \N__52445\ : std_logic;
signal \N__52442\ : std_logic;
signal \N__52439\ : std_logic;
signal \N__52432\ : std_logic;
signal \N__52427\ : std_logic;
signal \N__52426\ : std_logic;
signal \N__52425\ : std_logic;
signal \N__52424\ : std_logic;
signal \N__52423\ : std_logic;
signal \N__52422\ : std_logic;
signal \N__52421\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52419\ : std_logic;
signal \N__52418\ : std_logic;
signal \N__52417\ : std_logic;
signal \N__52416\ : std_logic;
signal \N__52413\ : std_logic;
signal \N__52408\ : std_logic;
signal \N__52405\ : std_logic;
signal \N__52402\ : std_logic;
signal \N__52401\ : std_logic;
signal \N__52400\ : std_logic;
signal \N__52397\ : std_logic;
signal \N__52394\ : std_logic;
signal \N__52389\ : std_logic;
signal \N__52388\ : std_logic;
signal \N__52387\ : std_logic;
signal \N__52384\ : std_logic;
signal \N__52379\ : std_logic;
signal \N__52376\ : std_logic;
signal \N__52375\ : std_logic;
signal \N__52374\ : std_logic;
signal \N__52373\ : std_logic;
signal \N__52372\ : std_logic;
signal \N__52371\ : std_logic;
signal \N__52370\ : std_logic;
signal \N__52369\ : std_logic;
signal \N__52368\ : std_logic;
signal \N__52367\ : std_logic;
signal \N__52366\ : std_logic;
signal \N__52365\ : std_logic;
signal \N__52364\ : std_logic;
signal \N__52363\ : std_logic;
signal \N__52362\ : std_logic;
signal \N__52361\ : std_logic;
signal \N__52358\ : std_logic;
signal \N__52355\ : std_logic;
signal \N__52352\ : std_logic;
signal \N__52347\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52339\ : std_logic;
signal \N__52332\ : std_logic;
signal \N__52329\ : std_logic;
signal \N__52326\ : std_logic;
signal \N__52323\ : std_logic;
signal \N__52320\ : std_logic;
signal \N__52307\ : std_logic;
signal \N__52304\ : std_logic;
signal \N__52291\ : std_logic;
signal \N__52284\ : std_logic;
signal \N__52275\ : std_logic;
signal \N__52268\ : std_logic;
signal \N__52253\ : std_logic;
signal \N__52250\ : std_logic;
signal \N__52247\ : std_logic;
signal \N__52244\ : std_logic;
signal \N__52241\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52239\ : std_logic;
signal \N__52238\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52236\ : std_logic;
signal \N__52235\ : std_logic;
signal \N__52234\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52230\ : std_logic;
signal \N__52227\ : std_logic;
signal \N__52224\ : std_logic;
signal \N__52223\ : std_logic;
signal \N__52222\ : std_logic;
signal \N__52221\ : std_logic;
signal \N__52216\ : std_logic;
signal \N__52215\ : std_logic;
signal \N__52214\ : std_logic;
signal \N__52213\ : std_logic;
signal \N__52212\ : std_logic;
signal \N__52211\ : std_logic;
signal \N__52210\ : std_logic;
signal \N__52209\ : std_logic;
signal \N__52208\ : std_logic;
signal \N__52207\ : std_logic;
signal \N__52206\ : std_logic;
signal \N__52205\ : std_logic;
signal \N__52204\ : std_logic;
signal \N__52201\ : std_logic;
signal \N__52198\ : std_logic;
signal \N__52197\ : std_logic;
signal \N__52196\ : std_logic;
signal \N__52191\ : std_logic;
signal \N__52190\ : std_logic;
signal \N__52189\ : std_logic;
signal \N__52188\ : std_logic;
signal \N__52187\ : std_logic;
signal \N__52184\ : std_logic;
signal \N__52181\ : std_logic;
signal \N__52178\ : std_logic;
signal \N__52173\ : std_logic;
signal \N__52170\ : std_logic;
signal \N__52167\ : std_logic;
signal \N__52154\ : std_logic;
signal \N__52141\ : std_logic;
signal \N__52136\ : std_logic;
signal \N__52131\ : std_logic;
signal \N__52128\ : std_logic;
signal \N__52125\ : std_logic;
signal \N__52122\ : std_logic;
signal \N__52117\ : std_logic;
signal \N__52112\ : std_logic;
signal \N__52109\ : std_logic;
signal \N__52106\ : std_logic;
signal \N__52095\ : std_logic;
signal \N__52090\ : std_logic;
signal \N__52073\ : std_logic;
signal \N__52072\ : std_logic;
signal \N__52069\ : std_logic;
signal \N__52068\ : std_logic;
signal \N__52065\ : std_logic;
signal \N__52062\ : std_logic;
signal \N__52059\ : std_logic;
signal \N__52058\ : std_logic;
signal \N__52055\ : std_logic;
signal \N__52050\ : std_logic;
signal \N__52047\ : std_logic;
signal \N__52044\ : std_logic;
signal \N__52039\ : std_logic;
signal \N__52036\ : std_logic;
signal \N__52033\ : std_logic;
signal \N__52030\ : std_logic;
signal \N__52027\ : std_logic;
signal \N__52022\ : std_logic;
signal \N__52021\ : std_logic;
signal \N__52016\ : std_logic;
signal \N__52013\ : std_logic;
signal \N__52010\ : std_logic;
signal \N__52009\ : std_logic;
signal \N__52006\ : std_logic;
signal \N__52003\ : std_logic;
signal \N__52000\ : std_logic;
signal \N__51995\ : std_logic;
signal \N__51992\ : std_logic;
signal \N__51989\ : std_logic;
signal \N__51986\ : std_logic;
signal \N__51985\ : std_logic;
signal \N__51980\ : std_logic;
signal \N__51977\ : std_logic;
signal \N__51974\ : std_logic;
signal \N__51973\ : std_logic;
signal \N__51968\ : std_logic;
signal \N__51965\ : std_logic;
signal \N__51962\ : std_logic;
signal \N__51959\ : std_logic;
signal \N__51956\ : std_logic;
signal \N__51953\ : std_logic;
signal \N__51950\ : std_logic;
signal \N__51949\ : std_logic;
signal \N__51946\ : std_logic;
signal \N__51943\ : std_logic;
signal \N__51938\ : std_logic;
signal \N__51935\ : std_logic;
signal \N__51932\ : std_logic;
signal \N__51929\ : std_logic;
signal \N__51928\ : std_logic;
signal \N__51925\ : std_logic;
signal \N__51922\ : std_logic;
signal \N__51919\ : std_logic;
signal \N__51916\ : std_logic;
signal \N__51911\ : std_logic;
signal \N__51908\ : std_logic;
signal \N__51907\ : std_logic;
signal \N__51902\ : std_logic;
signal \N__51899\ : std_logic;
signal \N__51896\ : std_logic;
signal \N__51895\ : std_logic;
signal \N__51890\ : std_logic;
signal \N__51887\ : std_logic;
signal \N__51884\ : std_logic;
signal \N__51881\ : std_logic;
signal \N__51878\ : std_logic;
signal \N__51877\ : std_logic;
signal \N__51874\ : std_logic;
signal \N__51871\ : std_logic;
signal \N__51866\ : std_logic;
signal \N__51863\ : std_logic;
signal \N__51860\ : std_logic;
signal \N__51859\ : std_logic;
signal \N__51856\ : std_logic;
signal \N__51853\ : std_logic;
signal \N__51850\ : std_logic;
signal \N__51847\ : std_logic;
signal \N__51842\ : std_logic;
signal \N__51841\ : std_logic;
signal \N__51836\ : std_logic;
signal \N__51833\ : std_logic;
signal \N__51830\ : std_logic;
signal \N__51829\ : std_logic;
signal \N__51824\ : std_logic;
signal \N__51821\ : std_logic;
signal \N__51818\ : std_logic;
signal \N__51815\ : std_logic;
signal \N__51814\ : std_logic;
signal \N__51813\ : std_logic;
signal \N__51810\ : std_logic;
signal \N__51805\ : std_logic;
signal \N__51804\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51798\ : std_logic;
signal \N__51795\ : std_logic;
signal \N__51790\ : std_logic;
signal \N__51785\ : std_logic;
signal \N__51782\ : std_logic;
signal \N__51781\ : std_logic;
signal \N__51780\ : std_logic;
signal \N__51777\ : std_logic;
signal \N__51772\ : std_logic;
signal \N__51771\ : std_logic;
signal \N__51768\ : std_logic;
signal \N__51765\ : std_logic;
signal \N__51762\ : std_logic;
signal \N__51757\ : std_logic;
signal \N__51752\ : std_logic;
signal \N__51749\ : std_logic;
signal \N__51748\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51746\ : std_logic;
signal \N__51743\ : std_logic;
signal \N__51740\ : std_logic;
signal \N__51737\ : std_logic;
signal \N__51734\ : std_logic;
signal \N__51731\ : std_logic;
signal \N__51728\ : std_logic;
signal \N__51723\ : std_logic;
signal \N__51720\ : std_logic;
signal \N__51717\ : std_logic;
signal \N__51714\ : std_logic;
signal \N__51707\ : std_logic;
signal \N__51706\ : std_logic;
signal \N__51705\ : std_logic;
signal \N__51702\ : std_logic;
signal \N__51699\ : std_logic;
signal \N__51696\ : std_logic;
signal \N__51693\ : std_logic;
signal \N__51690\ : std_logic;
signal \N__51689\ : std_logic;
signal \N__51684\ : std_logic;
signal \N__51681\ : std_logic;
signal \N__51678\ : std_logic;
signal \N__51675\ : std_logic;
signal \N__51668\ : std_logic;
signal \N__51665\ : std_logic;
signal \N__51664\ : std_logic;
signal \N__51661\ : std_logic;
signal \N__51660\ : std_logic;
signal \N__51657\ : std_logic;
signal \N__51656\ : std_logic;
signal \N__51653\ : std_logic;
signal \N__51650\ : std_logic;
signal \N__51647\ : std_logic;
signal \N__51644\ : std_logic;
signal \N__51641\ : std_logic;
signal \N__51638\ : std_logic;
signal \N__51629\ : std_logic;
signal \N__51628\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51622\ : std_logic;
signal \N__51619\ : std_logic;
signal \N__51618\ : std_logic;
signal \N__51615\ : std_logic;
signal \N__51612\ : std_logic;
signal \N__51609\ : std_logic;
signal \N__51602\ : std_logic;
signal \N__51599\ : std_logic;
signal \N__51596\ : std_logic;
signal \N__51595\ : std_logic;
signal \N__51594\ : std_logic;
signal \N__51593\ : std_logic;
signal \N__51590\ : std_logic;
signal \N__51587\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51579\ : std_logic;
signal \N__51576\ : std_logic;
signal \N__51569\ : std_logic;
signal \N__51566\ : std_logic;
signal \N__51563\ : std_logic;
signal \N__51562\ : std_logic;
signal \N__51559\ : std_logic;
signal \N__51556\ : std_logic;
signal \N__51555\ : std_logic;
signal \N__51552\ : std_logic;
signal \N__51549\ : std_logic;
signal \N__51546\ : std_logic;
signal \N__51539\ : std_logic;
signal \N__51536\ : std_logic;
signal \N__51535\ : std_logic;
signal \N__51534\ : std_logic;
signal \N__51531\ : std_logic;
signal \N__51528\ : std_logic;
signal \N__51525\ : std_logic;
signal \N__51522\ : std_logic;
signal \N__51519\ : std_logic;
signal \N__51518\ : std_logic;
signal \N__51515\ : std_logic;
signal \N__51510\ : std_logic;
signal \N__51507\ : std_logic;
signal \N__51500\ : std_logic;
signal \N__51497\ : std_logic;
signal \N__51496\ : std_logic;
signal \N__51495\ : std_logic;
signal \N__51492\ : std_logic;
signal \N__51489\ : std_logic;
signal \N__51486\ : std_logic;
signal \N__51483\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51475\ : std_logic;
signal \N__51474\ : std_logic;
signal \N__51471\ : std_logic;
signal \N__51468\ : std_logic;
signal \N__51465\ : std_logic;
signal \N__51458\ : std_logic;
signal \N__51455\ : std_logic;
signal \N__51452\ : std_logic;
signal \N__51449\ : std_logic;
signal \N__51446\ : std_logic;
signal \N__51443\ : std_logic;
signal \N__51440\ : std_logic;
signal \N__51437\ : std_logic;
signal \N__51436\ : std_logic;
signal \N__51433\ : std_logic;
signal \N__51432\ : std_logic;
signal \N__51431\ : std_logic;
signal \N__51428\ : std_logic;
signal \N__51425\ : std_logic;
signal \N__51422\ : std_logic;
signal \N__51419\ : std_logic;
signal \N__51416\ : std_logic;
signal \N__51407\ : std_logic;
signal \N__51404\ : std_logic;
signal \N__51401\ : std_logic;
signal \N__51398\ : std_logic;
signal \N__51395\ : std_logic;
signal \N__51392\ : std_logic;
signal \N__51389\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51379\ : std_logic;
signal \N__51378\ : std_logic;
signal \N__51377\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51368\ : std_logic;
signal \N__51365\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51359\ : std_logic;
signal \N__51356\ : std_logic;
signal \N__51353\ : std_logic;
signal \N__51346\ : std_logic;
signal \N__51341\ : std_logic;
signal \N__51338\ : std_logic;
signal \N__51335\ : std_logic;
signal \N__51332\ : std_logic;
signal \N__51331\ : std_logic;
signal \N__51328\ : std_logic;
signal \N__51325\ : std_logic;
signal \N__51324\ : std_logic;
signal \N__51321\ : std_logic;
signal \N__51316\ : std_logic;
signal \N__51315\ : std_logic;
signal \N__51312\ : std_logic;
signal \N__51309\ : std_logic;
signal \N__51306\ : std_logic;
signal \N__51301\ : std_logic;
signal \N__51298\ : std_logic;
signal \N__51293\ : std_logic;
signal \N__51290\ : std_logic;
signal \N__51287\ : std_logic;
signal \N__51284\ : std_logic;
signal \N__51281\ : std_logic;
signal \N__51280\ : std_logic;
signal \N__51277\ : std_logic;
signal \N__51276\ : std_logic;
signal \N__51275\ : std_logic;
signal \N__51272\ : std_logic;
signal \N__51269\ : std_logic;
signal \N__51264\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51254\ : std_logic;
signal \N__51251\ : std_logic;
signal \N__51248\ : std_logic;
signal \N__51245\ : std_logic;
signal \N__51242\ : std_logic;
signal \N__51239\ : std_logic;
signal \N__51236\ : std_logic;
signal \N__51233\ : std_logic;
signal \N__51232\ : std_logic;
signal \N__51231\ : std_logic;
signal \N__51230\ : std_logic;
signal \N__51227\ : std_logic;
signal \N__51224\ : std_logic;
signal \N__51219\ : std_logic;
signal \N__51212\ : std_logic;
signal \N__51209\ : std_logic;
signal \N__51206\ : std_logic;
signal \N__51203\ : std_logic;
signal \N__51200\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51196\ : std_logic;
signal \N__51193\ : std_logic;
signal \N__51190\ : std_logic;
signal \N__51189\ : std_logic;
signal \N__51188\ : std_logic;
signal \N__51185\ : std_logic;
signal \N__51182\ : std_logic;
signal \N__51179\ : std_logic;
signal \N__51176\ : std_logic;
signal \N__51167\ : std_logic;
signal \N__51164\ : std_logic;
signal \N__51161\ : std_logic;
signal \N__51158\ : std_logic;
signal \N__51155\ : std_logic;
signal \N__51152\ : std_logic;
signal \N__51149\ : std_logic;
signal \N__51148\ : std_logic;
signal \N__51145\ : std_logic;
signal \N__51142\ : std_logic;
signal \N__51141\ : std_logic;
signal \N__51140\ : std_logic;
signal \N__51137\ : std_logic;
signal \N__51134\ : std_logic;
signal \N__51131\ : std_logic;
signal \N__51128\ : std_logic;
signal \N__51119\ : std_logic;
signal \N__51116\ : std_logic;
signal \N__51113\ : std_logic;
signal \N__51110\ : std_logic;
signal \N__51107\ : std_logic;
signal \N__51104\ : std_logic;
signal \N__51101\ : std_logic;
signal \N__51100\ : std_logic;
signal \N__51097\ : std_logic;
signal \N__51096\ : std_logic;
signal \N__51093\ : std_logic;
signal \N__51092\ : std_logic;
signal \N__51089\ : std_logic;
signal \N__51086\ : std_logic;
signal \N__51081\ : std_logic;
signal \N__51074\ : std_logic;
signal \N__51071\ : std_logic;
signal \N__51070\ : std_logic;
signal \N__51067\ : std_logic;
signal \N__51064\ : std_logic;
signal \N__51063\ : std_logic;
signal \N__51062\ : std_logic;
signal \N__51059\ : std_logic;
signal \N__51056\ : std_logic;
signal \N__51053\ : std_logic;
signal \N__51050\ : std_logic;
signal \N__51041\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51035\ : std_logic;
signal \N__51032\ : std_logic;
signal \N__51029\ : std_logic;
signal \N__51026\ : std_logic;
signal \N__51023\ : std_logic;
signal \N__51020\ : std_logic;
signal \N__51017\ : std_logic;
signal \N__51014\ : std_logic;
signal \N__51011\ : std_logic;
signal \N__51008\ : std_logic;
signal \N__51005\ : std_logic;
signal \N__51002\ : std_logic;
signal \N__50999\ : std_logic;
signal \N__50996\ : std_logic;
signal \N__50993\ : std_logic;
signal \N__50990\ : std_logic;
signal \N__50987\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50981\ : std_logic;
signal \N__50978\ : std_logic;
signal \N__50975\ : std_logic;
signal \N__50972\ : std_logic;
signal \N__50969\ : std_logic;
signal \N__50966\ : std_logic;
signal \N__50963\ : std_logic;
signal \N__50960\ : std_logic;
signal \N__50957\ : std_logic;
signal \N__50954\ : std_logic;
signal \N__50951\ : std_logic;
signal \N__50950\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50946\ : std_logic;
signal \N__50945\ : std_logic;
signal \N__50940\ : std_logic;
signal \N__50937\ : std_logic;
signal \N__50934\ : std_logic;
signal \N__50931\ : std_logic;
signal \N__50924\ : std_logic;
signal \N__50921\ : std_logic;
signal \N__50918\ : std_logic;
signal \N__50915\ : std_logic;
signal \N__50912\ : std_logic;
signal \N__50909\ : std_logic;
signal \N__50906\ : std_logic;
signal \N__50905\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50903\ : std_logic;
signal \N__50900\ : std_logic;
signal \N__50897\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50889\ : std_logic;
signal \N__50884\ : std_logic;
signal \N__50879\ : std_logic;
signal \N__50876\ : std_logic;
signal \N__50873\ : std_logic;
signal \N__50870\ : std_logic;
signal \N__50867\ : std_logic;
signal \N__50864\ : std_logic;
signal \N__50861\ : std_logic;
signal \N__50858\ : std_logic;
signal \N__50855\ : std_logic;
signal \N__50852\ : std_logic;
signal \N__50849\ : std_logic;
signal \N__50848\ : std_logic;
signal \N__50845\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50840\ : std_logic;
signal \N__50837\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50829\ : std_logic;
signal \N__50826\ : std_logic;
signal \N__50823\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50813\ : std_logic;
signal \N__50810\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50804\ : std_logic;
signal \N__50801\ : std_logic;
signal \N__50798\ : std_logic;
signal \N__50795\ : std_logic;
signal \N__50794\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50787\ : std_logic;
signal \N__50786\ : std_logic;
signal \N__50783\ : std_logic;
signal \N__50780\ : std_logic;
signal \N__50777\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50765\ : std_logic;
signal \N__50762\ : std_logic;
signal \N__50759\ : std_logic;
signal \N__50756\ : std_logic;
signal \N__50753\ : std_logic;
signal \N__50750\ : std_logic;
signal \N__50749\ : std_logic;
signal \N__50748\ : std_logic;
signal \N__50747\ : std_logic;
signal \N__50744\ : std_logic;
signal \N__50741\ : std_logic;
signal \N__50736\ : std_logic;
signal \N__50731\ : std_logic;
signal \N__50728\ : std_logic;
signal \N__50725\ : std_logic;
signal \N__50720\ : std_logic;
signal \N__50717\ : std_logic;
signal \N__50714\ : std_logic;
signal \N__50711\ : std_logic;
signal \N__50708\ : std_logic;
signal \N__50705\ : std_logic;
signal \N__50702\ : std_logic;
signal \N__50699\ : std_logic;
signal \N__50696\ : std_logic;
signal \N__50693\ : std_logic;
signal \N__50692\ : std_logic;
signal \N__50689\ : std_logic;
signal \N__50686\ : std_logic;
signal \N__50685\ : std_logic;
signal \N__50682\ : std_logic;
signal \N__50681\ : std_logic;
signal \N__50678\ : std_logic;
signal \N__50675\ : std_logic;
signal \N__50672\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50664\ : std_logic;
signal \N__50661\ : std_logic;
signal \N__50658\ : std_logic;
signal \N__50655\ : std_logic;
signal \N__50648\ : std_logic;
signal \N__50645\ : std_logic;
signal \N__50642\ : std_logic;
signal \N__50639\ : std_logic;
signal \N__50636\ : std_logic;
signal \N__50633\ : std_logic;
signal \N__50630\ : std_logic;
signal \N__50629\ : std_logic;
signal \N__50626\ : std_logic;
signal \N__50623\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50619\ : std_logic;
signal \N__50618\ : std_logic;
signal \N__50615\ : std_logic;
signal \N__50612\ : std_logic;
signal \N__50609\ : std_logic;
signal \N__50606\ : std_logic;
signal \N__50603\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50591\ : std_logic;
signal \N__50588\ : std_logic;
signal \N__50585\ : std_logic;
signal \N__50582\ : std_logic;
signal \N__50579\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50572\ : std_logic;
signal \N__50571\ : std_logic;
signal \N__50570\ : std_logic;
signal \N__50565\ : std_logic;
signal \N__50562\ : std_logic;
signal \N__50559\ : std_logic;
signal \N__50556\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50540\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50534\ : std_logic;
signal \N__50531\ : std_logic;
signal \N__50528\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50522\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50511\ : std_logic;
signal \N__50508\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50492\ : std_logic;
signal \N__50489\ : std_logic;
signal \N__50486\ : std_logic;
signal \N__50483\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50471\ : std_logic;
signal \N__50468\ : std_logic;
signal \N__50465\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50459\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50450\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50444\ : std_logic;
signal \N__50441\ : std_logic;
signal \N__50438\ : std_logic;
signal \N__50435\ : std_logic;
signal \N__50432\ : std_logic;
signal \N__50429\ : std_logic;
signal \N__50426\ : std_logic;
signal \N__50423\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50414\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50399\ : std_logic;
signal \N__50396\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50360\ : std_logic;
signal \N__50357\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50350\ : std_logic;
signal \N__50347\ : std_logic;
signal \N__50344\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50258\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50216\ : std_logic;
signal \N__50213\ : std_logic;
signal \N__50210\ : std_logic;
signal \N__50207\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50203\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50194\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50186\ : std_logic;
signal \N__50185\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50176\ : std_logic;
signal \N__50171\ : std_logic;
signal \N__50168\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50164\ : std_logic;
signal \N__50159\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50155\ : std_logic;
signal \N__50152\ : std_logic;
signal \N__50149\ : std_logic;
signal \N__50146\ : std_logic;
signal \N__50141\ : std_logic;
signal \N__50138\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50136\ : std_logic;
signal \N__50135\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50127\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50125\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50121\ : std_logic;
signal \N__50120\ : std_logic;
signal \N__50119\ : std_logic;
signal \N__50118\ : std_logic;
signal \N__50117\ : std_logic;
signal \N__50112\ : std_logic;
signal \N__50111\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50104\ : std_logic;
signal \N__50103\ : std_logic;
signal \N__50102\ : std_logic;
signal \N__50101\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50099\ : std_logic;
signal \N__50098\ : std_logic;
signal \N__50097\ : std_logic;
signal \N__50096\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50091\ : std_logic;
signal \N__50090\ : std_logic;
signal \N__50089\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50087\ : std_logic;
signal \N__50086\ : std_logic;
signal \N__50085\ : std_logic;
signal \N__50084\ : std_logic;
signal \N__50083\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50081\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50065\ : std_logic;
signal \N__50060\ : std_logic;
signal \N__50059\ : std_logic;
signal \N__50050\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50046\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50025\ : std_logic;
signal \N__50022\ : std_logic;
signal \N__50021\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49997\ : std_logic;
signal \N__49996\ : std_logic;
signal \N__49995\ : std_logic;
signal \N__49994\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49992\ : std_logic;
signal \N__49991\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49989\ : std_logic;
signal \N__49988\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49985\ : std_logic;
signal \N__49982\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49980\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49973\ : std_logic;
signal \N__49970\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49951\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49945\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49937\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49935\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49912\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49804\ : std_logic;
signal \N__49801\ : std_logic;
signal \N__49796\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49769\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49766\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49761\ : std_logic;
signal \N__49760\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49757\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49751\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49728\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49724\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49716\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49713\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49708\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49705\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49667\ : std_logic;
signal \N__49662\ : std_logic;
signal \N__49651\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49649\ : std_logic;
signal \N__49640\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49635\ : std_logic;
signal \N__49634\ : std_logic;
signal \N__49631\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49625\ : std_logic;
signal \N__49624\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49622\ : std_logic;
signal \N__49621\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49619\ : std_logic;
signal \N__49618\ : std_logic;
signal \N__49617\ : std_logic;
signal \N__49616\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49614\ : std_logic;
signal \N__49613\ : std_logic;
signal \N__49612\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49606\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49592\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49572\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49563\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49560\ : std_logic;
signal \N__49559\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49557\ : std_logic;
signal \N__49556\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49553\ : std_logic;
signal \N__49552\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49550\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49547\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49544\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49541\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49535\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49511\ : std_logic;
signal \N__49510\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49508\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49502\ : std_logic;
signal \N__49501\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49492\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49487\ : std_logic;
signal \N__49484\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49463\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49421\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49409\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49399\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49358\ : std_logic;
signal \N__49355\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49347\ : std_logic;
signal \N__49346\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49339\ : std_logic;
signal \N__49338\ : std_logic;
signal \N__49335\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49330\ : std_logic;
signal \N__49327\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49322\ : std_logic;
signal \N__49319\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49315\ : std_logic;
signal \N__49314\ : std_logic;
signal \N__49301\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49287\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49277\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49234\ : std_logic;
signal \N__49217\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49157\ : std_logic;
signal \N__49154\ : std_logic;
signal \N__49151\ : std_logic;
signal \N__49148\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49118\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49097\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49085\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49072\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49062\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49052\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49036\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49032\ : std_logic;
signal \N__49031\ : std_logic;
signal \N__49028\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49010\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48995\ : std_logic;
signal \N__48992\ : std_logic;
signal \N__48989\ : std_logic;
signal \N__48986\ : std_logic;
signal \N__48983\ : std_logic;
signal \N__48982\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48965\ : std_logic;
signal \N__48964\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48947\ : std_logic;
signal \N__48944\ : std_logic;
signal \N__48941\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48923\ : std_logic;
signal \N__48920\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48905\ : std_logic;
signal \N__48902\ : std_logic;
signal \N__48899\ : std_logic;
signal \N__48896\ : std_logic;
signal \N__48893\ : std_logic;
signal \N__48890\ : std_logic;
signal \N__48887\ : std_logic;
signal \N__48884\ : std_logic;
signal \N__48881\ : std_logic;
signal \N__48878\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48850\ : std_logic;
signal \N__48849\ : std_logic;
signal \N__48842\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48827\ : std_logic;
signal \N__48824\ : std_logic;
signal \N__48821\ : std_logic;
signal \N__48818\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48794\ : std_logic;
signal \N__48793\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48772\ : std_logic;
signal \N__48771\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48747\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48744\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48726\ : std_logic;
signal \N__48725\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48690\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48644\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48605\ : std_logic;
signal \N__48602\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48593\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48584\ : std_logic;
signal \N__48581\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48560\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48521\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48515\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48506\ : std_logic;
signal \N__48503\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48491\ : std_logic;
signal \N__48488\ : std_logic;
signal \N__48485\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48476\ : std_logic;
signal \N__48473\ : std_logic;
signal \N__48470\ : std_logic;
signal \N__48467\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48455\ : std_logic;
signal \N__48452\ : std_logic;
signal \N__48449\ : std_logic;
signal \N__48446\ : std_logic;
signal \N__48443\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48434\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48428\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48398\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48380\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48374\ : std_logic;
signal \N__48371\ : std_logic;
signal \N__48368\ : std_logic;
signal \N__48365\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48359\ : std_logic;
signal \N__48356\ : std_logic;
signal \N__48353\ : std_logic;
signal \N__48350\ : std_logic;
signal \N__48347\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48320\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48302\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48281\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48245\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48230\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48218\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48209\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48200\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48116\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48107\ : std_logic;
signal \N__48104\ : std_logic;
signal \N__48101\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48083\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48077\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48071\ : std_logic;
signal \N__48068\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48062\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48053\ : std_logic;
signal \N__48050\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48044\ : std_logic;
signal \N__48041\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48035\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48008\ : std_logic;
signal \N__48005\ : std_logic;
signal \N__48002\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47975\ : std_logic;
signal \N__47972\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47966\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47942\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47936\ : std_logic;
signal \N__47933\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47717\ : std_logic;
signal \N__47714\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47525\ : std_logic;
signal \N__47522\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47513\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47504\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47459\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47441\ : std_logic;
signal \N__47438\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47417\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47303\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47219\ : std_logic;
signal \N__47216\ : std_logic;
signal \N__47213\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47207\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47198\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47186\ : std_logic;
signal \N__47183\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47177\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47171\ : std_logic;
signal \N__47168\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47159\ : std_logic;
signal \N__47156\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47129\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47114\ : std_logic;
signal \N__47111\ : std_logic;
signal \N__47108\ : std_logic;
signal \N__47105\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46952\ : std_logic;
signal \N__46949\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46838\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46721\ : std_logic;
signal \N__46718\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46685\ : std_logic;
signal \N__46682\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46592\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46577\ : std_logic;
signal \N__46574\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46556\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46499\ : std_logic;
signal \N__46496\ : std_logic;
signal \N__46493\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46472\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46451\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46436\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46430\ : std_logic;
signal \N__46427\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46421\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46400\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46337\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46313\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46286\ : std_logic;
signal \N__46283\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46262\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46244\ : std_logic;
signal \N__46241\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46226\ : std_logic;
signal \N__46223\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46187\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46088\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46073\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46006\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45973\ : std_logic;
signal \N__45970\ : std_logic;
signal \N__45967\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45921\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45901\ : std_logic;
signal \N__45898\ : std_logic;
signal \N__45895\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45828\ : std_logic;
signal \N__45823\ : std_logic;
signal \N__45820\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45808\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45776\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45772\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45761\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45754\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45709\ : std_logic;
signal \N__45706\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45679\ : std_logic;
signal \N__45676\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45652\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45518\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45421\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45395\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45328\ : std_logic;
signal \N__45319\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45217\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45171\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45160\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45062\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44809\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44780\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44747\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44743\ : std_logic;
signal \N__44740\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44690\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44686\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44680\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44630\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44521\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44284\ : std_logic;
signal \N__44281\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44192\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44101\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44024\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44011\ : std_logic;
signal \N__44008\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43999\ : std_logic;
signal \N__43996\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43918\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43868\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43631\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43624\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43537\ : std_logic;
signal \N__43534\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43394\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43247\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43214\ : std_logic;
signal \N__43211\ : std_logic;
signal \N__43208\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43181\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43172\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42911\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42719\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42685\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42596\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42553\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42343\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42211\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42107\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41977\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41966\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41909\ : std_logic;
signal \N__41906\ : std_logic;
signal \N__41903\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41870\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41528\ : std_logic;
signal \N__41525\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41483\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41459\ : std_logic;
signal \N__41456\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41450\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41411\ : std_logic;
signal \N__41408\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41300\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41273\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41165\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41134\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41110\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40823\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40780\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40682\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40646\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40581\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40568\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40560\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40286\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40219\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40055\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39956\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39871\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39672\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39487\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39481\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38063\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \pwm_generator_inst.O_0_1\ : std_logic;
signal \pwm_generator_inst.O_0_0\ : std_logic;
signal \pwm_generator_inst.O_0_5\ : std_logic;
signal \pwm_generator_inst.O_0_3\ : std_logic;
signal \pwm_generator_inst.O_0_4\ : std_logic;
signal \pwm_generator_inst.O_0_2\ : std_logic;
signal \pwm_generator_inst.O_0_6\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_0\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_8\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.O_11\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_11\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_15\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_19\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_20\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_21\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_22\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_23\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_24\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_25\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_20\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_22\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_21\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_15\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_15\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_23\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_8\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_25\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPFZ0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_15\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal \bfn_1_20_0_\ : std_logic;
signal \pwm_generator_inst.O_0_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CCZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_0_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DCZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_0_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI77ECZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.O_0_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FCZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.O_0_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGCZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.O_0_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHCZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.O_0_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFICZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FOZ0\ : std_logic;
signal \bfn_1_21_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDIZ0Z8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9_c_RNISHKZ0Z8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10_c_RNI59GZ0Z7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DIZ0Z7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HKZ0Z7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLMZ0Z7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPOZ0Z7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQZ0Z7\ : std_logic;
signal \bfn_1_22_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1TZ0Z7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFDZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNOZ0\ : std_logic;
signal \N_112_i_i\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_18\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_0_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_7\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_8_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_25\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_7_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_5_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_23\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_23\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_24\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_6_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_24\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_26\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSONZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_axb_16Z0Z_1_cascade_\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_1_15\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_25\ : std_logic;
signal un8_start_stop : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \bfn_3_12_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_3_13_0_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_1_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_19\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRROZ0\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_19\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_20\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_2_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_3_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_21\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_4_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_22\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0\ : std_logic;
signal \pwm_generator_inst.N_179_i\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_3_15_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.N_180_i\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.N_181_i\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.N_182_i\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.N_183_i\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.N_184_i\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.N_185_i\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.N_186_i\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.N_187_i\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_3_16_0_\ : std_logic;
signal \pwm_generator_inst.N_188_i\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_start_0\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst2.start_flagZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_0_sqmuxa\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_7\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_16\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_24\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_i_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0_g\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_0\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_8\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_30\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.measured_delay_tr_i_31\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_1 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_2 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_3 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_4 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_5 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_6 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_7 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_8 : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_9 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_10 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_11 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_12 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_13 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_14 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_15 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_16 : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_17 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_18 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_19 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_27 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_7\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_15\ : std_logic;
signal \bfn_8_22_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_23\ : std_logic;
signal \bfn_8_23_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0_g\ : std_logic;
signal s4_phy_c : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.state_ns_0_0_1\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_start_0\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal start_stop_c : std_logic;
signal \phase_controller_inst1.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst1.state_ns_0_0_1_cascade_\ : std_logic;
signal \phase_controller_inst1.start_flagZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIDC91B_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \elapsed_time_ns_1_RNIED91B_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_28 : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_0\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ1Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_8\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_30\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_24 : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_25 : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt26\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_26 : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_i_0\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal s3_phy_c : std_logic;
signal \bfn_10_2_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_7\ : std_logic;
signal \bfn_10_3_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_15\ : std_logic;
signal \bfn_10_4_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_23\ : std_logic;
signal \bfn_10_5_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_i_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_26\ : std_logic;
signal il_min_comp1_c : std_logic;
signal il_max_comp1_c : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \pwm_generator_inst.un3_threshold_iZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_20 : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_21 : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_22 : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_23 : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt20\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_0\ : std_logic;
signal \bfn_11_4_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_8\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_30\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_0\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ1Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_8\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_15\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_30\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_0\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_8\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_15\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_24\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \bfn_11_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_11_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.measured_delay_hc_i_31\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_1 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_5 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_8 : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_9 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_11 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_12 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_13 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_14 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_15 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_20 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_21 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_22 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_23 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_24 : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_26 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_27 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_4 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_4\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_2 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_2\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_6 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_6\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_19 : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_3 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_3\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_7 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_7\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_10 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_10\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_25 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_167_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt16\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_16 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_17 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt18\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_18 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_i_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_12_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_168_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ : std_logic;
signal \bfn_12_23_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ : std_logic;
signal \bfn_12_24_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\ : std_logic;
signal \GB_BUFFER_red_c_g_THRU_CO\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_28 : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt30\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_8\ : std_logic;
signal \bfn_13_21_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0\ : std_logic;
signal \bfn_13_22_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_CO\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13\ : std_logic;
signal \elapsed_time_ns_1_RNIDV2T9_0_1\ : std_logic;
signal \elapsed_time_ns_1_RNIE03T9_0_2\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.N_163_i_g\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_15\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_23\ : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \bfn_16_13_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\ : std_logic;
signal \bfn_16_14_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_17\ : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_9\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_3\ : std_logic;
signal \current_shift_inst.control_input_axb_0_cascade_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \bfn_17_3_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \bfn_17_4_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \bfn_17_5_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \bfn_17_6_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_165_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_17_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_166_i\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_8\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_16\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.N_1619_i\ : std_logic;
signal \current_shift_inst.control_input_1\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.control_input_axb_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.control_input_axb_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\ : std_logic;
signal \current_shift_inst.control_input_cry_13\ : std_logic;
signal \current_shift_inst.control_input_axb_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\ : std_logic;
signal \current_shift_inst.control_input_cry_14\ : std_logic;
signal \current_shift_inst.control_input_cry_15\ : std_logic;
signal \current_shift_inst.control_input_axb_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\ : std_logic;
signal \bfn_17_21_0_\ : std_logic;
signal \current_shift_inst.control_input_axb_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\ : std_logic;
signal \current_shift_inst.control_input_cry_16\ : std_logic;
signal \current_shift_inst.control_input_axb_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\ : std_logic;
signal \current_shift_inst.control_input_cry_17\ : std_logic;
signal \current_shift_inst.control_input_axb_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\ : std_logic;
signal \current_shift_inst.control_input_cry_18\ : std_logic;
signal \current_shift_inst.control_input_axb_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\ : std_logic;
signal \current_shift_inst.control_input_cry_19\ : std_logic;
signal \current_shift_inst.control_input_axb_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\ : std_logic;
signal \current_shift_inst.control_input_cry_20\ : std_logic;
signal \current_shift_inst.control_input_axb_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\ : std_logic;
signal \current_shift_inst.control_input_cry_21\ : std_logic;
signal \current_shift_inst.control_input_axb_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\ : std_logic;
signal \current_shift_inst.control_input_cry_22\ : std_logic;
signal \current_shift_inst.control_input_cry_23\ : std_logic;
signal \current_shift_inst.control_input_axb_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\ : std_logic;
signal \bfn_17_22_0_\ : std_logic;
signal \current_shift_inst.control_input_axb_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\ : std_logic;
signal \current_shift_inst.control_input_cry_24\ : std_logic;
signal \current_shift_inst.control_input_axb_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\ : std_logic;
signal \current_shift_inst.control_input_cry_25\ : std_logic;
signal \current_shift_inst.control_input_axb_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\ : std_logic;
signal \current_shift_inst.control_input_cry_26\ : std_logic;
signal \current_shift_inst.control_input_axb_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\ : std_logic;
signal \current_shift_inst.control_input_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\ : std_logic;
signal \current_shift_inst.control_input_cry_28\ : std_logic;
signal \current_shift_inst.control_input_cry_29\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.control_input_axb_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator\ : std_logic;
signal \bfn_17_23_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_9\ : std_logic;
signal \bfn_17_24_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_17\ : std_logic;
signal \bfn_17_25_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \bfn_17_26_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \current_shift_inst.timer_s1.N_164_i\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\ : std_logic;
signal state_3 : std_logic;
signal s1_phy_c : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.N_163_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \bfn_18_23_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \bfn_18_24_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \bfn_18_25_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \bfn_18_26_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_77_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal \current_shift_inst.PI_CTRL.N_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\ : std_logic;
signal pwm_duty_input_10 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal pwm_duty_input_8 : std_logic;
signal pwm_duty_input_3 : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal pwm_duty_input_1 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_94\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_120\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\ : std_logic_vector(31 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    pwm_output <= pwm_output_wire;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ <= \N__40358\&\N__40283\&\N__43367\&\N__40259\&\N__40481\&\N__40454\&\N__43391\&\N__43346\&\N__43502\&\N__40310\&\N__40337\&\N__40235\&\N__43475\&\N__40160\&\N__43325\&\N__43442\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__42347\&'0'&\N__42346\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_A_wire\ <= '0'&\N__52734\&\N__52737\&\N__52735\&\N__52738\&\N__52736\&\N__52853\&\N__52970\&\N__52667\&\N__53063\&\N__53009\&\N__52952\&\N__52964\&\N__52913\&\N__52934\&\N__52958\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__42763\&'0'&\N__42762\;
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(15);
    \pwm_generator_inst.O_0_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(14);
    \pwm_generator_inst.O_0_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(13);
    \pwm_generator_inst.O_0_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(12);
    \pwm_generator_inst.O_0_11\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(11);
    \pwm_generator_inst.O_0_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(10);
    \pwm_generator_inst.O_0_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(9);
    \pwm_generator_inst.O_0_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(8);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(7);
    \pwm_generator_inst.O_0_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(6);
    \pwm_generator_inst.O_0_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(5);
    \pwm_generator_inst.O_0_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(4);
    \pwm_generator_inst.O_0_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(3);
    \pwm_generator_inst.O_0_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(2);
    \pwm_generator_inst.O_0_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(1);
    \pwm_generator_inst.O_0_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_A_wire\ <= '0'&\N__22769\&\N__22805\&\N__22844\&\N__29846\&\N__21662\&\N__21746\&\N__21701\&\N__21722\&\N__21683\&\N__21788\&\N__21767\&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&\N__42481\&\N__42488\&\N__42484\&\N__42487\&\N__42482\&'0'&'0'&\N__42486\&\N__42483\&\N__42485\;
    \pwm_generator_inst.un5_threshold_1_26\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(26);
    \pwm_generator_inst.un5_threshold_1_25\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(25);
    \pwm_generator_inst.un5_threshold_1_24\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(24);
    \pwm_generator_inst.un5_threshold_1_23\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(23);
    \pwm_generator_inst.un5_threshold_1_22\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(22);
    \pwm_generator_inst.un5_threshold_1_21\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(21);
    \pwm_generator_inst.un5_threshold_1_20\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(20);
    \pwm_generator_inst.un5_threshold_1_19\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(19);
    \pwm_generator_inst.un5_threshold_1_18\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(18);
    \pwm_generator_inst.un5_threshold_1_17\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(17);
    \pwm_generator_inst.un5_threshold_1_16\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(16);
    \pwm_generator_inst.un5_threshold_1_15\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(12);
    \pwm_generator_inst.O_11\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_A_wire\ <= \N__52796\&\N__52788\&\N__52795\&\N__52787\&\N__52794\&\N__52786\&\N__52793\&\N__52785\&\N__52791\&\N__52783\&\N__52790\&\N__52784\&\N__52792\&\N__52782\&\N__52789\&\N__52781\;
    \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__42099\&'0'&\N__42098\;
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(0);
    \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_A_wire\ <= '0'&\N__23075\&\N__22874\&\N__22889\&\N__22904\&\N__22919\&\N__22934\&\N__22949\&\N__22964\&\N__22979\&\N__22994\&\N__22619\&\N__22634\&\N__22667\&\N__22703\&\N__22733\;
    \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&\N__41997\&\N__42004\&\N__42000\&\N__42003\&\N__41998\&'0'&'0'&\N__42002\&\N__41999\&\N__42001\;
    \pwm_generator_inst.un5_threshold_2_1_16\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(16);
    \pwm_generator_inst.un5_threshold_2_1_15\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(15);
    \pwm_generator_inst.un5_threshold_2_14\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(14);
    \pwm_generator_inst.un5_threshold_2_13\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(13);
    \pwm_generator_inst.un5_threshold_2_12\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(12);
    \pwm_generator_inst.un5_threshold_2_11\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(11);
    \pwm_generator_inst.un5_threshold_2_10\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(10);
    \pwm_generator_inst.un5_threshold_2_9\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(9);
    \pwm_generator_inst.un5_threshold_2_8\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(8);
    \pwm_generator_inst.un5_threshold_2_7\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(7);
    \pwm_generator_inst.un5_threshold_2_6\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(6);
    \pwm_generator_inst.un5_threshold_2_5\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(5);
    \pwm_generator_inst.un5_threshold_2_4\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(4);
    \pwm_generator_inst.un5_threshold_2_3\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(3);
    \pwm_generator_inst.un5_threshold_2_2\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(2);
    \pwm_generator_inst.un5_threshold_2_1\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(1);
    \pwm_generator_inst.un5_threshold_2_0\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(0);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ <= '0'&\N__50375\&\N__43526\&\N__50309\&\N__50258\&\N__50213\&\N__50357\&\N__50282\&\N__48923\&\N__48965\&\N__43421\&\N__48947\&\N__50333\&\N__50237\&\N__48989\&\N__53891\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__42607\&'0'&\N__42606\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(19);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(18);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(17);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(16);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.un1_integrator\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__23306\,
            RESETB => \N__35876\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42212\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__42345\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42704\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__42761\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42489\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__42480\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_A_wire\,
            C => \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_C_wire\,
            B => \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42091\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__42097\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\
        );

    \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42019\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__41996\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_A_wire\,
            C => \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_C_wire\,
            B => \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42211\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__42605\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__54405\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54407\,
            DIN => \N__54406\,
            DOUT => \N__54405\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54407\,
            PADOUT => \N__54406\,
            PADIN => \N__54405\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54396\,
            DIN => \N__54395\,
            DOUT => \N__54394\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54396\,
            PADOUT => \N__54395\,
            PADIN => \N__54394\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24023\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54387\,
            DIN => \N__54386\,
            DOUT => \N__54385\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54387\,
            PADOUT => \N__54386\,
            PADIN => \N__54385\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54378\,
            DIN => \N__54377\,
            DOUT => \N__54376\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54378\,
            PADOUT => \N__54377\,
            PADIN => \N__54376\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__49097\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54369\,
            DIN => \N__54368\,
            DOUT => \N__54367\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54369\,
            PADOUT => \N__54368\,
            PADIN => \N__54367\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26609\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54360\,
            DIN => \N__54359\,
            DOUT => \N__54358\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54360\,
            PADOUT => \N__54359\,
            PADIN => \N__54358\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54351\,
            DIN => \N__54350\,
            DOUT => \N__54349\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54351\,
            PADOUT => \N__54350\,
            PADIN => \N__54349\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28670\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54342\,
            DIN => \N__54341\,
            DOUT => \N__54340\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54342\,
            PADOUT => \N__54341\,
            PADIN => \N__54340\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54333\,
            DIN => \N__54332\,
            DOUT => \N__54331\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54333\,
            PADOUT => \N__54332\,
            PADIN => \N__54331\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54324\,
            DIN => \N__54323\,
            DOUT => \N__54322\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54324\,
            PADOUT => \N__54323\,
            PADIN => \N__54322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54315\,
            DIN => \N__54314\,
            DOUT => \N__54313\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54315\,
            PADOUT => \N__54314\,
            PADIN => \N__54313\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__30698\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54306\,
            DIN => \N__54305\,
            DOUT => \N__54304\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54306\,
            PADOUT => \N__54305\,
            PADIN => \N__54304\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54297\,
            DIN => \N__54296\,
            DOUT => \N__54295\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54297\,
            PADOUT => \N__54296\,
            PADIN => \N__54295\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__12659\ : CascadeMux
    port map (
            O => \N__54278\,
            I => \N__54275\
        );

    \I__12658\ : InMux
    port map (
            O => \N__54275\,
            I => \N__54269\
        );

    \I__12657\ : InMux
    port map (
            O => \N__54274\,
            I => \N__54269\
        );

    \I__12656\ : LocalMux
    port map (
            O => \N__54269\,
            I => \N__54266\
        );

    \I__12655\ : Odrv4
    port map (
            O => \N__54266\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__12654\ : InMux
    port map (
            O => \N__54263\,
            I => \N__54252\
        );

    \I__12653\ : InMux
    port map (
            O => \N__54262\,
            I => \N__54252\
        );

    \I__12652\ : InMux
    port map (
            O => \N__54261\,
            I => \N__54252\
        );

    \I__12651\ : CascadeMux
    port map (
            O => \N__54260\,
            I => \N__54249\
        );

    \I__12650\ : InMux
    port map (
            O => \N__54259\,
            I => \N__54243\
        );

    \I__12649\ : LocalMux
    port map (
            O => \N__54252\,
            I => \N__54240\
        );

    \I__12648\ : InMux
    port map (
            O => \N__54249\,
            I => \N__54237\
        );

    \I__12647\ : InMux
    port map (
            O => \N__54248\,
            I => \N__54232\
        );

    \I__12646\ : InMux
    port map (
            O => \N__54247\,
            I => \N__54232\
        );

    \I__12645\ : InMux
    port map (
            O => \N__54246\,
            I => \N__54229\
        );

    \I__12644\ : LocalMux
    port map (
            O => \N__54243\,
            I => \N__54222\
        );

    \I__12643\ : Span4Mux_v
    port map (
            O => \N__54240\,
            I => \N__54222\
        );

    \I__12642\ : LocalMux
    port map (
            O => \N__54237\,
            I => \N__54222\
        );

    \I__12641\ : LocalMux
    port map (
            O => \N__54232\,
            I => \N__54217\
        );

    \I__12640\ : LocalMux
    port map (
            O => \N__54229\,
            I => \N__54217\
        );

    \I__12639\ : Span4Mux_h
    port map (
            O => \N__54222\,
            I => \N__54214\
        );

    \I__12638\ : Span4Mux_s2_h
    port map (
            O => \N__54217\,
            I => \N__54211\
        );

    \I__12637\ : Span4Mux_v
    port map (
            O => \N__54214\,
            I => \N__54208\
        );

    \I__12636\ : Span4Mux_v
    port map (
            O => \N__54211\,
            I => \N__54205\
        );

    \I__12635\ : Span4Mux_v
    port map (
            O => \N__54208\,
            I => \N__54202\
        );

    \I__12634\ : Span4Mux_v
    port map (
            O => \N__54205\,
            I => \N__54199\
        );

    \I__12633\ : Odrv4
    port map (
            O => \N__54202\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10\
        );

    \I__12632\ : Odrv4
    port map (
            O => \N__54199\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10\
        );

    \I__12631\ : CascadeMux
    port map (
            O => \N__54194\,
            I => \current_shift_inst.PI_CTRL.N_97_cascade_\
        );

    \I__12630\ : InMux
    port map (
            O => \N__54191\,
            I => \N__54187\
        );

    \I__12629\ : InMux
    port map (
            O => \N__54190\,
            I => \N__54184\
        );

    \I__12628\ : LocalMux
    port map (
            O => \N__54187\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__12627\ : LocalMux
    port map (
            O => \N__54184\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__12626\ : InMux
    port map (
            O => \N__54179\,
            I => \N__54170\
        );

    \I__12625\ : InMux
    port map (
            O => \N__54178\,
            I => \N__54170\
        );

    \I__12624\ : InMux
    port map (
            O => \N__54177\,
            I => \N__54170\
        );

    \I__12623\ : LocalMux
    port map (
            O => \N__54170\,
            I => \current_shift_inst.PI_CTRL.N_120\
        );

    \I__12622\ : InMux
    port map (
            O => \N__54167\,
            I => \N__54161\
        );

    \I__12621\ : InMux
    port map (
            O => \N__54166\,
            I => \N__54158\
        );

    \I__12620\ : InMux
    port map (
            O => \N__54165\,
            I => \N__54155\
        );

    \I__12619\ : InMux
    port map (
            O => \N__54164\,
            I => \N__54152\
        );

    \I__12618\ : LocalMux
    port map (
            O => \N__54161\,
            I => \N__54147\
        );

    \I__12617\ : LocalMux
    port map (
            O => \N__54158\,
            I => \N__54147\
        );

    \I__12616\ : LocalMux
    port map (
            O => \N__54155\,
            I => \N__54144\
        );

    \I__12615\ : LocalMux
    port map (
            O => \N__54152\,
            I => \N__54141\
        );

    \I__12614\ : Span4Mux_v
    port map (
            O => \N__54147\,
            I => \N__54138\
        );

    \I__12613\ : Span4Mux_v
    port map (
            O => \N__54144\,
            I => \N__54133\
        );

    \I__12612\ : Span4Mux_s2_h
    port map (
            O => \N__54141\,
            I => \N__54133\
        );

    \I__12611\ : Span4Mux_v
    port map (
            O => \N__54138\,
            I => \N__54130\
        );

    \I__12610\ : Span4Mux_v
    port map (
            O => \N__54133\,
            I => \N__54127\
        );

    \I__12609\ : Span4Mux_h
    port map (
            O => \N__54130\,
            I => \N__54124\
        );

    \I__12608\ : Span4Mux_h
    port map (
            O => \N__54127\,
            I => \N__54121\
        );

    \I__12607\ : Odrv4
    port map (
            O => \N__54124\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__12606\ : Odrv4
    port map (
            O => \N__54121\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__12605\ : InMux
    port map (
            O => \N__54116\,
            I => \N__54111\
        );

    \I__12604\ : InMux
    port map (
            O => \N__54115\,
            I => \N__54108\
        );

    \I__12603\ : InMux
    port map (
            O => \N__54114\,
            I => \N__54105\
        );

    \I__12602\ : LocalMux
    port map (
            O => \N__54111\,
            I => \N__54098\
        );

    \I__12601\ : LocalMux
    port map (
            O => \N__54108\,
            I => \N__54098\
        );

    \I__12600\ : LocalMux
    port map (
            O => \N__54105\,
            I => \N__54098\
        );

    \I__12599\ : Span12Mux_v
    port map (
            O => \N__54098\,
            I => \N__54095\
        );

    \I__12598\ : Odrv12
    port map (
            O => \N__54095\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__12597\ : InMux
    port map (
            O => \N__54092\,
            I => \N__54080\
        );

    \I__12596\ : InMux
    port map (
            O => \N__54091\,
            I => \N__54080\
        );

    \I__12595\ : InMux
    port map (
            O => \N__54090\,
            I => \N__54073\
        );

    \I__12594\ : InMux
    port map (
            O => \N__54089\,
            I => \N__54073\
        );

    \I__12593\ : InMux
    port map (
            O => \N__54088\,
            I => \N__54073\
        );

    \I__12592\ : InMux
    port map (
            O => \N__54087\,
            I => \N__54068\
        );

    \I__12591\ : InMux
    port map (
            O => \N__54086\,
            I => \N__54068\
        );

    \I__12590\ : InMux
    port map (
            O => \N__54085\,
            I => \N__54064\
        );

    \I__12589\ : LocalMux
    port map (
            O => \N__54080\,
            I => \N__54056\
        );

    \I__12588\ : LocalMux
    port map (
            O => \N__54073\,
            I => \N__54056\
        );

    \I__12587\ : LocalMux
    port map (
            O => \N__54068\,
            I => \N__54056\
        );

    \I__12586\ : InMux
    port map (
            O => \N__54067\,
            I => \N__54053\
        );

    \I__12585\ : LocalMux
    port map (
            O => \N__54064\,
            I => \N__54050\
        );

    \I__12584\ : InMux
    port map (
            O => \N__54063\,
            I => \N__54047\
        );

    \I__12583\ : Span4Mux_v
    port map (
            O => \N__54056\,
            I => \N__54042\
        );

    \I__12582\ : LocalMux
    port map (
            O => \N__54053\,
            I => \N__54042\
        );

    \I__12581\ : Span4Mux_v
    port map (
            O => \N__54050\,
            I => \N__54037\
        );

    \I__12580\ : LocalMux
    port map (
            O => \N__54047\,
            I => \N__54037\
        );

    \I__12579\ : Span4Mux_h
    port map (
            O => \N__54042\,
            I => \N__54034\
        );

    \I__12578\ : Span4Mux_v
    port map (
            O => \N__54037\,
            I => \N__54031\
        );

    \I__12577\ : Span4Mux_v
    port map (
            O => \N__54034\,
            I => \N__54028\
        );

    \I__12576\ : Span4Mux_v
    port map (
            O => \N__54031\,
            I => \N__54025\
        );

    \I__12575\ : Span4Mux_v
    port map (
            O => \N__54028\,
            I => \N__54022\
        );

    \I__12574\ : Span4Mux_h
    port map (
            O => \N__54025\,
            I => \N__54019\
        );

    \I__12573\ : Odrv4
    port map (
            O => \N__54022\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__12572\ : Odrv4
    port map (
            O => \N__54019\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__12571\ : InMux
    port map (
            O => \N__54014\,
            I => \N__54011\
        );

    \I__12570\ : LocalMux
    port map (
            O => \N__54011\,
            I => \N__54007\
        );

    \I__12569\ : InMux
    port map (
            O => \N__54010\,
            I => \N__54004\
        );

    \I__12568\ : Odrv4
    port map (
            O => \N__54007\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__12567\ : LocalMux
    port map (
            O => \N__54004\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__12566\ : CascadeMux
    port map (
            O => \N__53999\,
            I => \current_shift_inst.PI_CTRL.N_98_cascade_\
        );

    \I__12565\ : CascadeMux
    port map (
            O => \N__53996\,
            I => \N__53989\
        );

    \I__12564\ : CascadeMux
    port map (
            O => \N__53995\,
            I => \N__53986\
        );

    \I__12563\ : CascadeMux
    port map (
            O => \N__53994\,
            I => \N__53983\
        );

    \I__12562\ : InMux
    port map (
            O => \N__53993\,
            I => \N__53979\
        );

    \I__12561\ : InMux
    port map (
            O => \N__53992\,
            I => \N__53976\
        );

    \I__12560\ : InMux
    port map (
            O => \N__53989\,
            I => \N__53973\
        );

    \I__12559\ : InMux
    port map (
            O => \N__53986\,
            I => \N__53966\
        );

    \I__12558\ : InMux
    port map (
            O => \N__53983\,
            I => \N__53966\
        );

    \I__12557\ : InMux
    port map (
            O => \N__53982\,
            I => \N__53966\
        );

    \I__12556\ : LocalMux
    port map (
            O => \N__53979\,
            I => \N__53960\
        );

    \I__12555\ : LocalMux
    port map (
            O => \N__53976\,
            I => \N__53960\
        );

    \I__12554\ : LocalMux
    port map (
            O => \N__53973\,
            I => \N__53957\
        );

    \I__12553\ : LocalMux
    port map (
            O => \N__53966\,
            I => \N__53954\
        );

    \I__12552\ : InMux
    port map (
            O => \N__53965\,
            I => \N__53951\
        );

    \I__12551\ : Span4Mux_s2_h
    port map (
            O => \N__53960\,
            I => \N__53948\
        );

    \I__12550\ : Span4Mux_s2_h
    port map (
            O => \N__53957\,
            I => \N__53943\
        );

    \I__12549\ : Span4Mux_s2_h
    port map (
            O => \N__53954\,
            I => \N__53943\
        );

    \I__12548\ : LocalMux
    port map (
            O => \N__53951\,
            I => \N__53940\
        );

    \I__12547\ : Span4Mux_v
    port map (
            O => \N__53948\,
            I => \N__53937\
        );

    \I__12546\ : Span4Mux_v
    port map (
            O => \N__53943\,
            I => \N__53934\
        );

    \I__12545\ : Span4Mux_s2_h
    port map (
            O => \N__53940\,
            I => \N__53931\
        );

    \I__12544\ : Span4Mux_v
    port map (
            O => \N__53937\,
            I => \N__53928\
        );

    \I__12543\ : Span4Mux_v
    port map (
            O => \N__53934\,
            I => \N__53925\
        );

    \I__12542\ : Span4Mux_v
    port map (
            O => \N__53931\,
            I => \N__53922\
        );

    \I__12541\ : Odrv4
    port map (
            O => \N__53928\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__12540\ : Odrv4
    port map (
            O => \N__53925\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__12539\ : Odrv4
    port map (
            O => \N__53922\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__12538\ : InMux
    port map (
            O => \N__53915\,
            I => \N__53912\
        );

    \I__12537\ : LocalMux
    port map (
            O => \N__53912\,
            I => \N__53908\
        );

    \I__12536\ : InMux
    port map (
            O => \N__53911\,
            I => \N__53905\
        );

    \I__12535\ : Odrv4
    port map (
            O => \N__53908\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__12534\ : LocalMux
    port map (
            O => \N__53905\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__12533\ : InMux
    port map (
            O => \N__53900\,
            I => \N__53897\
        );

    \I__12532\ : LocalMux
    port map (
            O => \N__53897\,
            I => \N__53894\
        );

    \I__12531\ : Odrv12
    port map (
            O => \N__53894\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__12530\ : InMux
    port map (
            O => \N__53891\,
            I => \N__53887\
        );

    \I__12529\ : InMux
    port map (
            O => \N__53890\,
            I => \N__53884\
        );

    \I__12528\ : LocalMux
    port map (
            O => \N__53887\,
            I => \N__53881\
        );

    \I__12527\ : LocalMux
    port map (
            O => \N__53884\,
            I => \N__53878\
        );

    \I__12526\ : Span4Mux_v
    port map (
            O => \N__53881\,
            I => \N__53875\
        );

    \I__12525\ : Span4Mux_h
    port map (
            O => \N__53878\,
            I => \N__53872\
        );

    \I__12524\ : Span4Mux_h
    port map (
            O => \N__53875\,
            I => \N__53869\
        );

    \I__12523\ : Span4Mux_h
    port map (
            O => \N__53872\,
            I => \N__53864\
        );

    \I__12522\ : Span4Mux_h
    port map (
            O => \N__53869\,
            I => \N__53864\
        );

    \I__12521\ : Odrv4
    port map (
            O => \N__53864\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__12520\ : InMux
    port map (
            O => \N__53861\,
            I => \N__53858\
        );

    \I__12519\ : LocalMux
    port map (
            O => \N__53858\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__12518\ : ClkMux
    port map (
            O => \N__53855\,
            I => \N__53468\
        );

    \I__12517\ : ClkMux
    port map (
            O => \N__53854\,
            I => \N__53468\
        );

    \I__12516\ : ClkMux
    port map (
            O => \N__53853\,
            I => \N__53468\
        );

    \I__12515\ : ClkMux
    port map (
            O => \N__53852\,
            I => \N__53468\
        );

    \I__12514\ : ClkMux
    port map (
            O => \N__53851\,
            I => \N__53468\
        );

    \I__12513\ : ClkMux
    port map (
            O => \N__53850\,
            I => \N__53468\
        );

    \I__12512\ : ClkMux
    port map (
            O => \N__53849\,
            I => \N__53468\
        );

    \I__12511\ : ClkMux
    port map (
            O => \N__53848\,
            I => \N__53468\
        );

    \I__12510\ : ClkMux
    port map (
            O => \N__53847\,
            I => \N__53468\
        );

    \I__12509\ : ClkMux
    port map (
            O => \N__53846\,
            I => \N__53468\
        );

    \I__12508\ : ClkMux
    port map (
            O => \N__53845\,
            I => \N__53468\
        );

    \I__12507\ : ClkMux
    port map (
            O => \N__53844\,
            I => \N__53468\
        );

    \I__12506\ : ClkMux
    port map (
            O => \N__53843\,
            I => \N__53468\
        );

    \I__12505\ : ClkMux
    port map (
            O => \N__53842\,
            I => \N__53468\
        );

    \I__12504\ : ClkMux
    port map (
            O => \N__53841\,
            I => \N__53468\
        );

    \I__12503\ : ClkMux
    port map (
            O => \N__53840\,
            I => \N__53468\
        );

    \I__12502\ : ClkMux
    port map (
            O => \N__53839\,
            I => \N__53468\
        );

    \I__12501\ : ClkMux
    port map (
            O => \N__53838\,
            I => \N__53468\
        );

    \I__12500\ : ClkMux
    port map (
            O => \N__53837\,
            I => \N__53468\
        );

    \I__12499\ : ClkMux
    port map (
            O => \N__53836\,
            I => \N__53468\
        );

    \I__12498\ : ClkMux
    port map (
            O => \N__53835\,
            I => \N__53468\
        );

    \I__12497\ : ClkMux
    port map (
            O => \N__53834\,
            I => \N__53468\
        );

    \I__12496\ : ClkMux
    port map (
            O => \N__53833\,
            I => \N__53468\
        );

    \I__12495\ : ClkMux
    port map (
            O => \N__53832\,
            I => \N__53468\
        );

    \I__12494\ : ClkMux
    port map (
            O => \N__53831\,
            I => \N__53468\
        );

    \I__12493\ : ClkMux
    port map (
            O => \N__53830\,
            I => \N__53468\
        );

    \I__12492\ : ClkMux
    port map (
            O => \N__53829\,
            I => \N__53468\
        );

    \I__12491\ : ClkMux
    port map (
            O => \N__53828\,
            I => \N__53468\
        );

    \I__12490\ : ClkMux
    port map (
            O => \N__53827\,
            I => \N__53468\
        );

    \I__12489\ : ClkMux
    port map (
            O => \N__53826\,
            I => \N__53468\
        );

    \I__12488\ : ClkMux
    port map (
            O => \N__53825\,
            I => \N__53468\
        );

    \I__12487\ : ClkMux
    port map (
            O => \N__53824\,
            I => \N__53468\
        );

    \I__12486\ : ClkMux
    port map (
            O => \N__53823\,
            I => \N__53468\
        );

    \I__12485\ : ClkMux
    port map (
            O => \N__53822\,
            I => \N__53468\
        );

    \I__12484\ : ClkMux
    port map (
            O => \N__53821\,
            I => \N__53468\
        );

    \I__12483\ : ClkMux
    port map (
            O => \N__53820\,
            I => \N__53468\
        );

    \I__12482\ : ClkMux
    port map (
            O => \N__53819\,
            I => \N__53468\
        );

    \I__12481\ : ClkMux
    port map (
            O => \N__53818\,
            I => \N__53468\
        );

    \I__12480\ : ClkMux
    port map (
            O => \N__53817\,
            I => \N__53468\
        );

    \I__12479\ : ClkMux
    port map (
            O => \N__53816\,
            I => \N__53468\
        );

    \I__12478\ : ClkMux
    port map (
            O => \N__53815\,
            I => \N__53468\
        );

    \I__12477\ : ClkMux
    port map (
            O => \N__53814\,
            I => \N__53468\
        );

    \I__12476\ : ClkMux
    port map (
            O => \N__53813\,
            I => \N__53468\
        );

    \I__12475\ : ClkMux
    port map (
            O => \N__53812\,
            I => \N__53468\
        );

    \I__12474\ : ClkMux
    port map (
            O => \N__53811\,
            I => \N__53468\
        );

    \I__12473\ : ClkMux
    port map (
            O => \N__53810\,
            I => \N__53468\
        );

    \I__12472\ : ClkMux
    port map (
            O => \N__53809\,
            I => \N__53468\
        );

    \I__12471\ : ClkMux
    port map (
            O => \N__53808\,
            I => \N__53468\
        );

    \I__12470\ : ClkMux
    port map (
            O => \N__53807\,
            I => \N__53468\
        );

    \I__12469\ : ClkMux
    port map (
            O => \N__53806\,
            I => \N__53468\
        );

    \I__12468\ : ClkMux
    port map (
            O => \N__53805\,
            I => \N__53468\
        );

    \I__12467\ : ClkMux
    port map (
            O => \N__53804\,
            I => \N__53468\
        );

    \I__12466\ : ClkMux
    port map (
            O => \N__53803\,
            I => \N__53468\
        );

    \I__12465\ : ClkMux
    port map (
            O => \N__53802\,
            I => \N__53468\
        );

    \I__12464\ : ClkMux
    port map (
            O => \N__53801\,
            I => \N__53468\
        );

    \I__12463\ : ClkMux
    port map (
            O => \N__53800\,
            I => \N__53468\
        );

    \I__12462\ : ClkMux
    port map (
            O => \N__53799\,
            I => \N__53468\
        );

    \I__12461\ : ClkMux
    port map (
            O => \N__53798\,
            I => \N__53468\
        );

    \I__12460\ : ClkMux
    port map (
            O => \N__53797\,
            I => \N__53468\
        );

    \I__12459\ : ClkMux
    port map (
            O => \N__53796\,
            I => \N__53468\
        );

    \I__12458\ : ClkMux
    port map (
            O => \N__53795\,
            I => \N__53468\
        );

    \I__12457\ : ClkMux
    port map (
            O => \N__53794\,
            I => \N__53468\
        );

    \I__12456\ : ClkMux
    port map (
            O => \N__53793\,
            I => \N__53468\
        );

    \I__12455\ : ClkMux
    port map (
            O => \N__53792\,
            I => \N__53468\
        );

    \I__12454\ : ClkMux
    port map (
            O => \N__53791\,
            I => \N__53468\
        );

    \I__12453\ : ClkMux
    port map (
            O => \N__53790\,
            I => \N__53468\
        );

    \I__12452\ : ClkMux
    port map (
            O => \N__53789\,
            I => \N__53468\
        );

    \I__12451\ : ClkMux
    port map (
            O => \N__53788\,
            I => \N__53468\
        );

    \I__12450\ : ClkMux
    port map (
            O => \N__53787\,
            I => \N__53468\
        );

    \I__12449\ : ClkMux
    port map (
            O => \N__53786\,
            I => \N__53468\
        );

    \I__12448\ : ClkMux
    port map (
            O => \N__53785\,
            I => \N__53468\
        );

    \I__12447\ : ClkMux
    port map (
            O => \N__53784\,
            I => \N__53468\
        );

    \I__12446\ : ClkMux
    port map (
            O => \N__53783\,
            I => \N__53468\
        );

    \I__12445\ : ClkMux
    port map (
            O => \N__53782\,
            I => \N__53468\
        );

    \I__12444\ : ClkMux
    port map (
            O => \N__53781\,
            I => \N__53468\
        );

    \I__12443\ : ClkMux
    port map (
            O => \N__53780\,
            I => \N__53468\
        );

    \I__12442\ : ClkMux
    port map (
            O => \N__53779\,
            I => \N__53468\
        );

    \I__12441\ : ClkMux
    port map (
            O => \N__53778\,
            I => \N__53468\
        );

    \I__12440\ : ClkMux
    port map (
            O => \N__53777\,
            I => \N__53468\
        );

    \I__12439\ : ClkMux
    port map (
            O => \N__53776\,
            I => \N__53468\
        );

    \I__12438\ : ClkMux
    port map (
            O => \N__53775\,
            I => \N__53468\
        );

    \I__12437\ : ClkMux
    port map (
            O => \N__53774\,
            I => \N__53468\
        );

    \I__12436\ : ClkMux
    port map (
            O => \N__53773\,
            I => \N__53468\
        );

    \I__12435\ : ClkMux
    port map (
            O => \N__53772\,
            I => \N__53468\
        );

    \I__12434\ : ClkMux
    port map (
            O => \N__53771\,
            I => \N__53468\
        );

    \I__12433\ : ClkMux
    port map (
            O => \N__53770\,
            I => \N__53468\
        );

    \I__12432\ : ClkMux
    port map (
            O => \N__53769\,
            I => \N__53468\
        );

    \I__12431\ : ClkMux
    port map (
            O => \N__53768\,
            I => \N__53468\
        );

    \I__12430\ : ClkMux
    port map (
            O => \N__53767\,
            I => \N__53468\
        );

    \I__12429\ : ClkMux
    port map (
            O => \N__53766\,
            I => \N__53468\
        );

    \I__12428\ : ClkMux
    port map (
            O => \N__53765\,
            I => \N__53468\
        );

    \I__12427\ : ClkMux
    port map (
            O => \N__53764\,
            I => \N__53468\
        );

    \I__12426\ : ClkMux
    port map (
            O => \N__53763\,
            I => \N__53468\
        );

    \I__12425\ : ClkMux
    port map (
            O => \N__53762\,
            I => \N__53468\
        );

    \I__12424\ : ClkMux
    port map (
            O => \N__53761\,
            I => \N__53468\
        );

    \I__12423\ : ClkMux
    port map (
            O => \N__53760\,
            I => \N__53468\
        );

    \I__12422\ : ClkMux
    port map (
            O => \N__53759\,
            I => \N__53468\
        );

    \I__12421\ : ClkMux
    port map (
            O => \N__53758\,
            I => \N__53468\
        );

    \I__12420\ : ClkMux
    port map (
            O => \N__53757\,
            I => \N__53468\
        );

    \I__12419\ : ClkMux
    port map (
            O => \N__53756\,
            I => \N__53468\
        );

    \I__12418\ : ClkMux
    port map (
            O => \N__53755\,
            I => \N__53468\
        );

    \I__12417\ : ClkMux
    port map (
            O => \N__53754\,
            I => \N__53468\
        );

    \I__12416\ : ClkMux
    port map (
            O => \N__53753\,
            I => \N__53468\
        );

    \I__12415\ : ClkMux
    port map (
            O => \N__53752\,
            I => \N__53468\
        );

    \I__12414\ : ClkMux
    port map (
            O => \N__53751\,
            I => \N__53468\
        );

    \I__12413\ : ClkMux
    port map (
            O => \N__53750\,
            I => \N__53468\
        );

    \I__12412\ : ClkMux
    port map (
            O => \N__53749\,
            I => \N__53468\
        );

    \I__12411\ : ClkMux
    port map (
            O => \N__53748\,
            I => \N__53468\
        );

    \I__12410\ : ClkMux
    port map (
            O => \N__53747\,
            I => \N__53468\
        );

    \I__12409\ : ClkMux
    port map (
            O => \N__53746\,
            I => \N__53468\
        );

    \I__12408\ : ClkMux
    port map (
            O => \N__53745\,
            I => \N__53468\
        );

    \I__12407\ : ClkMux
    port map (
            O => \N__53744\,
            I => \N__53468\
        );

    \I__12406\ : ClkMux
    port map (
            O => \N__53743\,
            I => \N__53468\
        );

    \I__12405\ : ClkMux
    port map (
            O => \N__53742\,
            I => \N__53468\
        );

    \I__12404\ : ClkMux
    port map (
            O => \N__53741\,
            I => \N__53468\
        );

    \I__12403\ : ClkMux
    port map (
            O => \N__53740\,
            I => \N__53468\
        );

    \I__12402\ : ClkMux
    port map (
            O => \N__53739\,
            I => \N__53468\
        );

    \I__12401\ : ClkMux
    port map (
            O => \N__53738\,
            I => \N__53468\
        );

    \I__12400\ : ClkMux
    port map (
            O => \N__53737\,
            I => \N__53468\
        );

    \I__12399\ : ClkMux
    port map (
            O => \N__53736\,
            I => \N__53468\
        );

    \I__12398\ : ClkMux
    port map (
            O => \N__53735\,
            I => \N__53468\
        );

    \I__12397\ : ClkMux
    port map (
            O => \N__53734\,
            I => \N__53468\
        );

    \I__12396\ : ClkMux
    port map (
            O => \N__53733\,
            I => \N__53468\
        );

    \I__12395\ : ClkMux
    port map (
            O => \N__53732\,
            I => \N__53468\
        );

    \I__12394\ : ClkMux
    port map (
            O => \N__53731\,
            I => \N__53468\
        );

    \I__12393\ : ClkMux
    port map (
            O => \N__53730\,
            I => \N__53468\
        );

    \I__12392\ : ClkMux
    port map (
            O => \N__53729\,
            I => \N__53468\
        );

    \I__12391\ : ClkMux
    port map (
            O => \N__53728\,
            I => \N__53468\
        );

    \I__12390\ : ClkMux
    port map (
            O => \N__53727\,
            I => \N__53468\
        );

    \I__12389\ : GlobalMux
    port map (
            O => \N__53468\,
            I => clk_100mhz_0
        );

    \I__12388\ : InMux
    port map (
            O => \N__53465\,
            I => \N__53455\
        );

    \I__12387\ : InMux
    port map (
            O => \N__53464\,
            I => \N__53452\
        );

    \I__12386\ : InMux
    port map (
            O => \N__53463\,
            I => \N__53449\
        );

    \I__12385\ : InMux
    port map (
            O => \N__53462\,
            I => \N__53446\
        );

    \I__12384\ : InMux
    port map (
            O => \N__53461\,
            I => \N__53443\
        );

    \I__12383\ : InMux
    port map (
            O => \N__53460\,
            I => \N__53440\
        );

    \I__12382\ : InMux
    port map (
            O => \N__53459\,
            I => \N__53437\
        );

    \I__12381\ : InMux
    port map (
            O => \N__53458\,
            I => \N__53434\
        );

    \I__12380\ : LocalMux
    port map (
            O => \N__53455\,
            I => \N__53431\
        );

    \I__12379\ : LocalMux
    port map (
            O => \N__53452\,
            I => \N__53428\
        );

    \I__12378\ : LocalMux
    port map (
            O => \N__53449\,
            I => \N__53425\
        );

    \I__12377\ : LocalMux
    port map (
            O => \N__53446\,
            I => \N__53419\
        );

    \I__12376\ : LocalMux
    port map (
            O => \N__53443\,
            I => \N__53397\
        );

    \I__12375\ : LocalMux
    port map (
            O => \N__53440\,
            I => \N__53359\
        );

    \I__12374\ : LocalMux
    port map (
            O => \N__53437\,
            I => \N__53351\
        );

    \I__12373\ : LocalMux
    port map (
            O => \N__53434\,
            I => \N__53332\
        );

    \I__12372\ : Glb2LocalMux
    port map (
            O => \N__53431\,
            I => \N__53099\
        );

    \I__12371\ : Glb2LocalMux
    port map (
            O => \N__53428\,
            I => \N__53099\
        );

    \I__12370\ : Glb2LocalMux
    port map (
            O => \N__53425\,
            I => \N__53099\
        );

    \I__12369\ : SRMux
    port map (
            O => \N__53424\,
            I => \N__53099\
        );

    \I__12368\ : SRMux
    port map (
            O => \N__53423\,
            I => \N__53099\
        );

    \I__12367\ : SRMux
    port map (
            O => \N__53422\,
            I => \N__53099\
        );

    \I__12366\ : Glb2LocalMux
    port map (
            O => \N__53419\,
            I => \N__53099\
        );

    \I__12365\ : SRMux
    port map (
            O => \N__53418\,
            I => \N__53099\
        );

    \I__12364\ : SRMux
    port map (
            O => \N__53417\,
            I => \N__53099\
        );

    \I__12363\ : SRMux
    port map (
            O => \N__53416\,
            I => \N__53099\
        );

    \I__12362\ : SRMux
    port map (
            O => \N__53415\,
            I => \N__53099\
        );

    \I__12361\ : SRMux
    port map (
            O => \N__53414\,
            I => \N__53099\
        );

    \I__12360\ : SRMux
    port map (
            O => \N__53413\,
            I => \N__53099\
        );

    \I__12359\ : SRMux
    port map (
            O => \N__53412\,
            I => \N__53099\
        );

    \I__12358\ : SRMux
    port map (
            O => \N__53411\,
            I => \N__53099\
        );

    \I__12357\ : SRMux
    port map (
            O => \N__53410\,
            I => \N__53099\
        );

    \I__12356\ : SRMux
    port map (
            O => \N__53409\,
            I => \N__53099\
        );

    \I__12355\ : SRMux
    port map (
            O => \N__53408\,
            I => \N__53099\
        );

    \I__12354\ : SRMux
    port map (
            O => \N__53407\,
            I => \N__53099\
        );

    \I__12353\ : SRMux
    port map (
            O => \N__53406\,
            I => \N__53099\
        );

    \I__12352\ : SRMux
    port map (
            O => \N__53405\,
            I => \N__53099\
        );

    \I__12351\ : SRMux
    port map (
            O => \N__53404\,
            I => \N__53099\
        );

    \I__12350\ : SRMux
    port map (
            O => \N__53403\,
            I => \N__53099\
        );

    \I__12349\ : SRMux
    port map (
            O => \N__53402\,
            I => \N__53099\
        );

    \I__12348\ : SRMux
    port map (
            O => \N__53401\,
            I => \N__53099\
        );

    \I__12347\ : SRMux
    port map (
            O => \N__53400\,
            I => \N__53099\
        );

    \I__12346\ : Glb2LocalMux
    port map (
            O => \N__53397\,
            I => \N__53099\
        );

    \I__12345\ : SRMux
    port map (
            O => \N__53396\,
            I => \N__53099\
        );

    \I__12344\ : SRMux
    port map (
            O => \N__53395\,
            I => \N__53099\
        );

    \I__12343\ : SRMux
    port map (
            O => \N__53394\,
            I => \N__53099\
        );

    \I__12342\ : SRMux
    port map (
            O => \N__53393\,
            I => \N__53099\
        );

    \I__12341\ : SRMux
    port map (
            O => \N__53392\,
            I => \N__53099\
        );

    \I__12340\ : SRMux
    port map (
            O => \N__53391\,
            I => \N__53099\
        );

    \I__12339\ : SRMux
    port map (
            O => \N__53390\,
            I => \N__53099\
        );

    \I__12338\ : SRMux
    port map (
            O => \N__53389\,
            I => \N__53099\
        );

    \I__12337\ : SRMux
    port map (
            O => \N__53388\,
            I => \N__53099\
        );

    \I__12336\ : SRMux
    port map (
            O => \N__53387\,
            I => \N__53099\
        );

    \I__12335\ : SRMux
    port map (
            O => \N__53386\,
            I => \N__53099\
        );

    \I__12334\ : SRMux
    port map (
            O => \N__53385\,
            I => \N__53099\
        );

    \I__12333\ : SRMux
    port map (
            O => \N__53384\,
            I => \N__53099\
        );

    \I__12332\ : SRMux
    port map (
            O => \N__53383\,
            I => \N__53099\
        );

    \I__12331\ : SRMux
    port map (
            O => \N__53382\,
            I => \N__53099\
        );

    \I__12330\ : SRMux
    port map (
            O => \N__53381\,
            I => \N__53099\
        );

    \I__12329\ : SRMux
    port map (
            O => \N__53380\,
            I => \N__53099\
        );

    \I__12328\ : SRMux
    port map (
            O => \N__53379\,
            I => \N__53099\
        );

    \I__12327\ : SRMux
    port map (
            O => \N__53378\,
            I => \N__53099\
        );

    \I__12326\ : SRMux
    port map (
            O => \N__53377\,
            I => \N__53099\
        );

    \I__12325\ : SRMux
    port map (
            O => \N__53376\,
            I => \N__53099\
        );

    \I__12324\ : SRMux
    port map (
            O => \N__53375\,
            I => \N__53099\
        );

    \I__12323\ : SRMux
    port map (
            O => \N__53374\,
            I => \N__53099\
        );

    \I__12322\ : SRMux
    port map (
            O => \N__53373\,
            I => \N__53099\
        );

    \I__12321\ : SRMux
    port map (
            O => \N__53372\,
            I => \N__53099\
        );

    \I__12320\ : SRMux
    port map (
            O => \N__53371\,
            I => \N__53099\
        );

    \I__12319\ : SRMux
    port map (
            O => \N__53370\,
            I => \N__53099\
        );

    \I__12318\ : SRMux
    port map (
            O => \N__53369\,
            I => \N__53099\
        );

    \I__12317\ : SRMux
    port map (
            O => \N__53368\,
            I => \N__53099\
        );

    \I__12316\ : SRMux
    port map (
            O => \N__53367\,
            I => \N__53099\
        );

    \I__12315\ : SRMux
    port map (
            O => \N__53366\,
            I => \N__53099\
        );

    \I__12314\ : SRMux
    port map (
            O => \N__53365\,
            I => \N__53099\
        );

    \I__12313\ : SRMux
    port map (
            O => \N__53364\,
            I => \N__53099\
        );

    \I__12312\ : SRMux
    port map (
            O => \N__53363\,
            I => \N__53099\
        );

    \I__12311\ : SRMux
    port map (
            O => \N__53362\,
            I => \N__53099\
        );

    \I__12310\ : Glb2LocalMux
    port map (
            O => \N__53359\,
            I => \N__53099\
        );

    \I__12309\ : SRMux
    port map (
            O => \N__53358\,
            I => \N__53099\
        );

    \I__12308\ : SRMux
    port map (
            O => \N__53357\,
            I => \N__53099\
        );

    \I__12307\ : SRMux
    port map (
            O => \N__53356\,
            I => \N__53099\
        );

    \I__12306\ : SRMux
    port map (
            O => \N__53355\,
            I => \N__53099\
        );

    \I__12305\ : SRMux
    port map (
            O => \N__53354\,
            I => \N__53099\
        );

    \I__12304\ : Glb2LocalMux
    port map (
            O => \N__53351\,
            I => \N__53099\
        );

    \I__12303\ : SRMux
    port map (
            O => \N__53350\,
            I => \N__53099\
        );

    \I__12302\ : SRMux
    port map (
            O => \N__53349\,
            I => \N__53099\
        );

    \I__12301\ : SRMux
    port map (
            O => \N__53348\,
            I => \N__53099\
        );

    \I__12300\ : SRMux
    port map (
            O => \N__53347\,
            I => \N__53099\
        );

    \I__12299\ : SRMux
    port map (
            O => \N__53346\,
            I => \N__53099\
        );

    \I__12298\ : SRMux
    port map (
            O => \N__53345\,
            I => \N__53099\
        );

    \I__12297\ : SRMux
    port map (
            O => \N__53344\,
            I => \N__53099\
        );

    \I__12296\ : SRMux
    port map (
            O => \N__53343\,
            I => \N__53099\
        );

    \I__12295\ : SRMux
    port map (
            O => \N__53342\,
            I => \N__53099\
        );

    \I__12294\ : SRMux
    port map (
            O => \N__53341\,
            I => \N__53099\
        );

    \I__12293\ : SRMux
    port map (
            O => \N__53340\,
            I => \N__53099\
        );

    \I__12292\ : SRMux
    port map (
            O => \N__53339\,
            I => \N__53099\
        );

    \I__12291\ : SRMux
    port map (
            O => \N__53338\,
            I => \N__53099\
        );

    \I__12290\ : SRMux
    port map (
            O => \N__53337\,
            I => \N__53099\
        );

    \I__12289\ : SRMux
    port map (
            O => \N__53336\,
            I => \N__53099\
        );

    \I__12288\ : SRMux
    port map (
            O => \N__53335\,
            I => \N__53099\
        );

    \I__12287\ : Glb2LocalMux
    port map (
            O => \N__53332\,
            I => \N__53099\
        );

    \I__12286\ : SRMux
    port map (
            O => \N__53331\,
            I => \N__53099\
        );

    \I__12285\ : SRMux
    port map (
            O => \N__53330\,
            I => \N__53099\
        );

    \I__12284\ : SRMux
    port map (
            O => \N__53329\,
            I => \N__53099\
        );

    \I__12283\ : SRMux
    port map (
            O => \N__53328\,
            I => \N__53099\
        );

    \I__12282\ : SRMux
    port map (
            O => \N__53327\,
            I => \N__53099\
        );

    \I__12281\ : SRMux
    port map (
            O => \N__53326\,
            I => \N__53099\
        );

    \I__12280\ : SRMux
    port map (
            O => \N__53325\,
            I => \N__53099\
        );

    \I__12279\ : SRMux
    port map (
            O => \N__53324\,
            I => \N__53099\
        );

    \I__12278\ : SRMux
    port map (
            O => \N__53323\,
            I => \N__53099\
        );

    \I__12277\ : SRMux
    port map (
            O => \N__53322\,
            I => \N__53099\
        );

    \I__12276\ : SRMux
    port map (
            O => \N__53321\,
            I => \N__53099\
        );

    \I__12275\ : SRMux
    port map (
            O => \N__53320\,
            I => \N__53099\
        );

    \I__12274\ : SRMux
    port map (
            O => \N__53319\,
            I => \N__53099\
        );

    \I__12273\ : SRMux
    port map (
            O => \N__53318\,
            I => \N__53099\
        );

    \I__12272\ : SRMux
    port map (
            O => \N__53317\,
            I => \N__53099\
        );

    \I__12271\ : SRMux
    port map (
            O => \N__53316\,
            I => \N__53099\
        );

    \I__12270\ : SRMux
    port map (
            O => \N__53315\,
            I => \N__53099\
        );

    \I__12269\ : SRMux
    port map (
            O => \N__53314\,
            I => \N__53099\
        );

    \I__12268\ : SRMux
    port map (
            O => \N__53313\,
            I => \N__53099\
        );

    \I__12267\ : SRMux
    port map (
            O => \N__53312\,
            I => \N__53099\
        );

    \I__12266\ : GlobalMux
    port map (
            O => \N__53099\,
            I => \N__53096\
        );

    \I__12265\ : gio2CtrlBuf
    port map (
            O => \N__53096\,
            I => red_c_g
        );

    \I__12264\ : InMux
    port map (
            O => \N__53093\,
            I => \N__53086\
        );

    \I__12263\ : InMux
    port map (
            O => \N__53092\,
            I => \N__53086\
        );

    \I__12262\ : InMux
    port map (
            O => \N__53091\,
            I => \N__53083\
        );

    \I__12261\ : LocalMux
    port map (
            O => \N__53086\,
            I => \N__53080\
        );

    \I__12260\ : LocalMux
    port map (
            O => \N__53083\,
            I => \N__53077\
        );

    \I__12259\ : Span4Mux_v
    port map (
            O => \N__53080\,
            I => \N__53074\
        );

    \I__12258\ : Span12Mux_s7_h
    port map (
            O => \N__53077\,
            I => \N__53071\
        );

    \I__12257\ : Span4Mux_h
    port map (
            O => \N__53074\,
            I => \N__53068\
        );

    \I__12256\ : Odrv12
    port map (
            O => \N__53071\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__12255\ : Odrv4
    port map (
            O => \N__53068\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__12254\ : InMux
    port map (
            O => \N__53063\,
            I => \N__53060\
        );

    \I__12253\ : LocalMux
    port map (
            O => \N__53060\,
            I => pwm_duty_input_6
        );

    \I__12252\ : CascadeMux
    port map (
            O => \N__53057\,
            I => \N__53053\
        );

    \I__12251\ : CascadeMux
    port map (
            O => \N__53056\,
            I => \N__53050\
        );

    \I__12250\ : InMux
    port map (
            O => \N__53053\,
            I => \N__53047\
        );

    \I__12249\ : InMux
    port map (
            O => \N__53050\,
            I => \N__53044\
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__53047\,
            I => \N__53040\
        );

    \I__12247\ : LocalMux
    port map (
            O => \N__53044\,
            I => \N__53037\
        );

    \I__12246\ : InMux
    port map (
            O => \N__53043\,
            I => \N__53034\
        );

    \I__12245\ : Span4Mux_v
    port map (
            O => \N__53040\,
            I => \N__53031\
        );

    \I__12244\ : Span4Mux_s2_h
    port map (
            O => \N__53037\,
            I => \N__53026\
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__53034\,
            I => \N__53026\
        );

    \I__12242\ : Span4Mux_v
    port map (
            O => \N__53031\,
            I => \N__53023\
        );

    \I__12241\ : Span4Mux_v
    port map (
            O => \N__53026\,
            I => \N__53020\
        );

    \I__12240\ : Span4Mux_h
    port map (
            O => \N__53023\,
            I => \N__53017\
        );

    \I__12239\ : Span4Mux_h
    port map (
            O => \N__53020\,
            I => \N__53014\
        );

    \I__12238\ : Odrv4
    port map (
            O => \N__53017\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__12237\ : Odrv4
    port map (
            O => \N__53014\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__12236\ : InMux
    port map (
            O => \N__53009\,
            I => \N__53006\
        );

    \I__12235\ : LocalMux
    port map (
            O => \N__53006\,
            I => pwm_duty_input_5
        );

    \I__12234\ : InMux
    port map (
            O => \N__53003\,
            I => \N__52999\
        );

    \I__12233\ : InMux
    port map (
            O => \N__53002\,
            I => \N__52996\
        );

    \I__12232\ : LocalMux
    port map (
            O => \N__52999\,
            I => \N__52993\
        );

    \I__12231\ : LocalMux
    port map (
            O => \N__52996\,
            I => \N__52990\
        );

    \I__12230\ : Span4Mux_v
    port map (
            O => \N__52993\,
            I => \N__52984\
        );

    \I__12229\ : Span4Mux_v
    port map (
            O => \N__52990\,
            I => \N__52984\
        );

    \I__12228\ : InMux
    port map (
            O => \N__52989\,
            I => \N__52981\
        );

    \I__12227\ : Sp12to4
    port map (
            O => \N__52984\,
            I => \N__52976\
        );

    \I__12226\ : LocalMux
    port map (
            O => \N__52981\,
            I => \N__52976\
        );

    \I__12225\ : Span12Mux_s7_h
    port map (
            O => \N__52976\,
            I => \N__52973\
        );

    \I__12224\ : Odrv12
    port map (
            O => \N__52973\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__12223\ : InMux
    port map (
            O => \N__52970\,
            I => \N__52967\
        );

    \I__12222\ : LocalMux
    port map (
            O => \N__52967\,
            I => pwm_duty_input_8
        );

    \I__12221\ : InMux
    port map (
            O => \N__52964\,
            I => \N__52961\
        );

    \I__12220\ : LocalMux
    port map (
            O => \N__52961\,
            I => pwm_duty_input_3
        );

    \I__12219\ : InMux
    port map (
            O => \N__52958\,
            I => \N__52955\
        );

    \I__12218\ : LocalMux
    port map (
            O => \N__52955\,
            I => pwm_duty_input_0
        );

    \I__12217\ : InMux
    port map (
            O => \N__52952\,
            I => \N__52949\
        );

    \I__12216\ : LocalMux
    port map (
            O => \N__52949\,
            I => pwm_duty_input_4
        );

    \I__12215\ : InMux
    port map (
            O => \N__52946\,
            I => \N__52943\
        );

    \I__12214\ : LocalMux
    port map (
            O => \N__52943\,
            I => \N__52940\
        );

    \I__12213\ : Span12Mux_s7_h
    port map (
            O => \N__52940\,
            I => \N__52937\
        );

    \I__12212\ : Odrv12
    port map (
            O => \N__52937\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__12211\ : InMux
    port map (
            O => \N__52934\,
            I => \N__52931\
        );

    \I__12210\ : LocalMux
    port map (
            O => \N__52931\,
            I => pwm_duty_input_1
        );

    \I__12209\ : InMux
    port map (
            O => \N__52928\,
            I => \N__52925\
        );

    \I__12208\ : LocalMux
    port map (
            O => \N__52925\,
            I => \N__52922\
        );

    \I__12207\ : Sp12to4
    port map (
            O => \N__52922\,
            I => \N__52919\
        );

    \I__12206\ : Span12Mux_v
    port map (
            O => \N__52919\,
            I => \N__52916\
        );

    \I__12205\ : Odrv12
    port map (
            O => \N__52916\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__12204\ : InMux
    port map (
            O => \N__52913\,
            I => \N__52910\
        );

    \I__12203\ : LocalMux
    port map (
            O => \N__52910\,
            I => pwm_duty_input_2
        );

    \I__12202\ : InMux
    port map (
            O => \N__52907\,
            I => \N__52904\
        );

    \I__12201\ : LocalMux
    port map (
            O => \N__52904\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__12200\ : InMux
    port map (
            O => \N__52901\,
            I => \N__52898\
        );

    \I__12199\ : LocalMux
    port map (
            O => \N__52898\,
            I => \N__52895\
        );

    \I__12198\ : Span4Mux_h
    port map (
            O => \N__52895\,
            I => \N__52892\
        );

    \I__12197\ : Odrv4
    port map (
            O => \N__52892\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__12196\ : InMux
    port map (
            O => \N__52889\,
            I => \N__52886\
        );

    \I__12195\ : LocalMux
    port map (
            O => \N__52886\,
            I => \N__52883\
        );

    \I__12194\ : Odrv4
    port map (
            O => \N__52883\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__12193\ : CascadeMux
    port map (
            O => \N__52880\,
            I => \N__52877\
        );

    \I__12192\ : InMux
    port map (
            O => \N__52877\,
            I => \N__52874\
        );

    \I__12191\ : LocalMux
    port map (
            O => \N__52874\,
            I => \N__52871\
        );

    \I__12190\ : Span4Mux_v
    port map (
            O => \N__52871\,
            I => \N__52868\
        );

    \I__12189\ : Odrv4
    port map (
            O => \N__52868\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__12188\ : InMux
    port map (
            O => \N__52865\,
            I => \N__52862\
        );

    \I__12187\ : LocalMux
    port map (
            O => \N__52862\,
            I => \N__52859\
        );

    \I__12186\ : Span4Mux_h
    port map (
            O => \N__52859\,
            I => \N__52856\
        );

    \I__12185\ : Odrv4
    port map (
            O => \N__52856\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__12184\ : InMux
    port map (
            O => \N__52853\,
            I => \N__52850\
        );

    \I__12183\ : LocalMux
    port map (
            O => \N__52850\,
            I => \N__52847\
        );

    \I__12182\ : Span4Mux_s1_h
    port map (
            O => \N__52847\,
            I => \N__52844\
        );

    \I__12181\ : Odrv4
    port map (
            O => \N__52844\,
            I => pwm_duty_input_9
        );

    \I__12180\ : CascadeMux
    port map (
            O => \N__52841\,
            I => \current_shift_inst.PI_CTRL.N_31_cascade_\
        );

    \I__12179\ : CascadeMux
    port map (
            O => \N__52838\,
            I => \N__52835\
        );

    \I__12178\ : InMux
    port map (
            O => \N__52835\,
            I => \N__52832\
        );

    \I__12177\ : LocalMux
    port map (
            O => \N__52832\,
            I => \N__52827\
        );

    \I__12176\ : InMux
    port map (
            O => \N__52831\,
            I => \N__52824\
        );

    \I__12175\ : InMux
    port map (
            O => \N__52830\,
            I => \N__52821\
        );

    \I__12174\ : Span4Mux_v
    port map (
            O => \N__52827\,
            I => \N__52814\
        );

    \I__12173\ : LocalMux
    port map (
            O => \N__52824\,
            I => \N__52814\
        );

    \I__12172\ : LocalMux
    port map (
            O => \N__52821\,
            I => \N__52814\
        );

    \I__12171\ : Span4Mux_v
    port map (
            O => \N__52814\,
            I => \N__52811\
        );

    \I__12170\ : Span4Mux_h
    port map (
            O => \N__52811\,
            I => \N__52808\
        );

    \I__12169\ : Odrv4
    port map (
            O => \N__52808\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__12168\ : CascadeMux
    port map (
            O => \N__52805\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\
        );

    \I__12167\ : InMux
    port map (
            O => \N__52802\,
            I => \N__52799\
        );

    \I__12166\ : LocalMux
    port map (
            O => \N__52799\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\
        );

    \I__12165\ : InMux
    port map (
            O => \N__52796\,
            I => \N__52764\
        );

    \I__12164\ : InMux
    port map (
            O => \N__52795\,
            I => \N__52764\
        );

    \I__12163\ : InMux
    port map (
            O => \N__52794\,
            I => \N__52764\
        );

    \I__12162\ : InMux
    port map (
            O => \N__52793\,
            I => \N__52764\
        );

    \I__12161\ : InMux
    port map (
            O => \N__52792\,
            I => \N__52764\
        );

    \I__12160\ : InMux
    port map (
            O => \N__52791\,
            I => \N__52764\
        );

    \I__12159\ : InMux
    port map (
            O => \N__52790\,
            I => \N__52764\
        );

    \I__12158\ : InMux
    port map (
            O => \N__52789\,
            I => \N__52764\
        );

    \I__12157\ : InMux
    port map (
            O => \N__52788\,
            I => \N__52747\
        );

    \I__12156\ : InMux
    port map (
            O => \N__52787\,
            I => \N__52747\
        );

    \I__12155\ : InMux
    port map (
            O => \N__52786\,
            I => \N__52747\
        );

    \I__12154\ : InMux
    port map (
            O => \N__52785\,
            I => \N__52747\
        );

    \I__12153\ : InMux
    port map (
            O => \N__52784\,
            I => \N__52747\
        );

    \I__12152\ : InMux
    port map (
            O => \N__52783\,
            I => \N__52747\
        );

    \I__12151\ : InMux
    port map (
            O => \N__52782\,
            I => \N__52747\
        );

    \I__12150\ : InMux
    port map (
            O => \N__52781\,
            I => \N__52747\
        );

    \I__12149\ : LocalMux
    port map (
            O => \N__52764\,
            I => \N__52742\
        );

    \I__12148\ : LocalMux
    port map (
            O => \N__52747\,
            I => \N__52742\
        );

    \I__12147\ : Span4Mux_v
    port map (
            O => \N__52742\,
            I => \N__52739\
        );

    \I__12146\ : Sp12to4
    port map (
            O => \N__52739\,
            I => \N__52731\
        );

    \I__12145\ : InMux
    port map (
            O => \N__52738\,
            I => \N__52726\
        );

    \I__12144\ : InMux
    port map (
            O => \N__52737\,
            I => \N__52726\
        );

    \I__12143\ : InMux
    port map (
            O => \N__52736\,
            I => \N__52719\
        );

    \I__12142\ : InMux
    port map (
            O => \N__52735\,
            I => \N__52719\
        );

    \I__12141\ : InMux
    port map (
            O => \N__52734\,
            I => \N__52719\
        );

    \I__12140\ : Span12Mux_s8_h
    port map (
            O => \N__52731\,
            I => \N__52716\
        );

    \I__12139\ : LocalMux
    port map (
            O => \N__52726\,
            I => \N__52711\
        );

    \I__12138\ : LocalMux
    port map (
            O => \N__52719\,
            I => \N__52711\
        );

    \I__12137\ : Span12Mux_h
    port map (
            O => \N__52716\,
            I => \N__52708\
        );

    \I__12136\ : Odrv4
    port map (
            O => \N__52711\,
            I => pwm_duty_input_10
        );

    \I__12135\ : Odrv12
    port map (
            O => \N__52708\,
            I => pwm_duty_input_10
        );

    \I__12134\ : InMux
    port map (
            O => \N__52703\,
            I => \N__52700\
        );

    \I__12133\ : LocalMux
    port map (
            O => \N__52700\,
            I => \N__52695\
        );

    \I__12132\ : InMux
    port map (
            O => \N__52699\,
            I => \N__52690\
        );

    \I__12131\ : InMux
    port map (
            O => \N__52698\,
            I => \N__52690\
        );

    \I__12130\ : Span4Mux_h
    port map (
            O => \N__52695\,
            I => \N__52687\
        );

    \I__12129\ : LocalMux
    port map (
            O => \N__52690\,
            I => \N__52684\
        );

    \I__12128\ : Span4Mux_v
    port map (
            O => \N__52687\,
            I => \N__52681\
        );

    \I__12127\ : Span4Mux_v
    port map (
            O => \N__52684\,
            I => \N__52678\
        );

    \I__12126\ : Span4Mux_v
    port map (
            O => \N__52681\,
            I => \N__52675\
        );

    \I__12125\ : Span4Mux_h
    port map (
            O => \N__52678\,
            I => \N__52672\
        );

    \I__12124\ : Odrv4
    port map (
            O => \N__52675\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__12123\ : Odrv4
    port map (
            O => \N__52672\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__12122\ : InMux
    port map (
            O => \N__52667\,
            I => \N__52664\
        );

    \I__12121\ : LocalMux
    port map (
            O => \N__52664\,
            I => \N__52661\
        );

    \I__12120\ : Odrv4
    port map (
            O => \N__52661\,
            I => pwm_duty_input_7
        );

    \I__12119\ : InMux
    port map (
            O => \N__52658\,
            I => \N__52655\
        );

    \I__12118\ : LocalMux
    port map (
            O => \N__52655\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__12117\ : CascadeMux
    port map (
            O => \N__52652\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\
        );

    \I__12116\ : InMux
    port map (
            O => \N__52649\,
            I => \N__52643\
        );

    \I__12115\ : InMux
    port map (
            O => \N__52648\,
            I => \N__52643\
        );

    \I__12114\ : LocalMux
    port map (
            O => \N__52643\,
            I => \N__52640\
        );

    \I__12113\ : Odrv4
    port map (
            O => \N__52640\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__12112\ : InMux
    port map (
            O => \N__52637\,
            I => \N__52634\
        );

    \I__12111\ : LocalMux
    port map (
            O => \N__52634\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__12110\ : InMux
    port map (
            O => \N__52631\,
            I => \N__52628\
        );

    \I__12109\ : LocalMux
    port map (
            O => \N__52628\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__12108\ : CascadeMux
    port map (
            O => \N__52625\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\
        );

    \I__12107\ : InMux
    port map (
            O => \N__52622\,
            I => \N__52618\
        );

    \I__12106\ : InMux
    port map (
            O => \N__52621\,
            I => \N__52615\
        );

    \I__12105\ : LocalMux
    port map (
            O => \N__52618\,
            I => \N__52612\
        );

    \I__12104\ : LocalMux
    port map (
            O => \N__52615\,
            I => \N__52609\
        );

    \I__12103\ : Span4Mux_h
    port map (
            O => \N__52612\,
            I => \N__52606\
        );

    \I__12102\ : Odrv4
    port map (
            O => \N__52609\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__12101\ : Odrv4
    port map (
            O => \N__52606\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__12100\ : InMux
    port map (
            O => \N__52601\,
            I => \N__52597\
        );

    \I__12099\ : InMux
    port map (
            O => \N__52600\,
            I => \N__52594\
        );

    \I__12098\ : LocalMux
    port map (
            O => \N__52597\,
            I => \N__52591\
        );

    \I__12097\ : LocalMux
    port map (
            O => \N__52594\,
            I => \N__52588\
        );

    \I__12096\ : Span4Mux_h
    port map (
            O => \N__52591\,
            I => \N__52585\
        );

    \I__12095\ : Odrv4
    port map (
            O => \N__52588\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__12094\ : Odrv4
    port map (
            O => \N__52585\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__12093\ : InMux
    port map (
            O => \N__52580\,
            I => \N__52576\
        );

    \I__12092\ : InMux
    port map (
            O => \N__52579\,
            I => \N__52573\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__52576\,
            I => \N__52570\
        );

    \I__12090\ : LocalMux
    port map (
            O => \N__52573\,
            I => \N__52567\
        );

    \I__12089\ : Span4Mux_h
    port map (
            O => \N__52570\,
            I => \N__52564\
        );

    \I__12088\ : Odrv4
    port map (
            O => \N__52567\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__12087\ : Odrv4
    port map (
            O => \N__52564\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__12086\ : CascadeMux
    port map (
            O => \N__52559\,
            I => \N__52555\
        );

    \I__12085\ : InMux
    port map (
            O => \N__52558\,
            I => \N__52550\
        );

    \I__12084\ : InMux
    port map (
            O => \N__52555\,
            I => \N__52550\
        );

    \I__12083\ : LocalMux
    port map (
            O => \N__52550\,
            I => \N__52547\
        );

    \I__12082\ : Odrv4
    port map (
            O => \N__52547\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__12081\ : InMux
    port map (
            O => \N__52544\,
            I => \N__52538\
        );

    \I__12080\ : InMux
    port map (
            O => \N__52543\,
            I => \N__52538\
        );

    \I__12079\ : LocalMux
    port map (
            O => \N__52538\,
            I => \N__52535\
        );

    \I__12078\ : Odrv4
    port map (
            O => \N__52535\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__12077\ : InMux
    port map (
            O => \N__52532\,
            I => \N__52526\
        );

    \I__12076\ : InMux
    port map (
            O => \N__52531\,
            I => \N__52526\
        );

    \I__12075\ : LocalMux
    port map (
            O => \N__52526\,
            I => \N__52523\
        );

    \I__12074\ : Odrv4
    port map (
            O => \N__52523\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__12073\ : InMux
    port map (
            O => \N__52520\,
            I => \N__52514\
        );

    \I__12072\ : InMux
    port map (
            O => \N__52519\,
            I => \N__52514\
        );

    \I__12071\ : LocalMux
    port map (
            O => \N__52514\,
            I => \N__52511\
        );

    \I__12070\ : Odrv4
    port map (
            O => \N__52511\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__12069\ : CascadeMux
    port map (
            O => \N__52508\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\
        );

    \I__12068\ : CascadeMux
    port map (
            O => \N__52505\,
            I => \N__52501\
        );

    \I__12067\ : InMux
    port map (
            O => \N__52504\,
            I => \N__52498\
        );

    \I__12066\ : InMux
    port map (
            O => \N__52501\,
            I => \N__52495\
        );

    \I__12065\ : LocalMux
    port map (
            O => \N__52498\,
            I => \N__52490\
        );

    \I__12064\ : LocalMux
    port map (
            O => \N__52495\,
            I => \N__52490\
        );

    \I__12063\ : Span4Mux_h
    port map (
            O => \N__52490\,
            I => \N__52487\
        );

    \I__12062\ : Odrv4
    port map (
            O => \N__52487\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__12061\ : InMux
    port map (
            O => \N__52484\,
            I => \N__52481\
        );

    \I__12060\ : LocalMux
    port map (
            O => \N__52481\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__12059\ : InMux
    port map (
            O => \N__52478\,
            I => \N__52475\
        );

    \I__12058\ : LocalMux
    port map (
            O => \N__52475\,
            I => \N__52472\
        );

    \I__12057\ : Span4Mux_h
    port map (
            O => \N__52472\,
            I => \N__52469\
        );

    \I__12056\ : Odrv4
    port map (
            O => \N__52469\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__12055\ : CascadeMux
    port map (
            O => \N__52466\,
            I => \N__52463\
        );

    \I__12054\ : InMux
    port map (
            O => \N__52463\,
            I => \N__52459\
        );

    \I__12053\ : InMux
    port map (
            O => \N__52462\,
            I => \N__52456\
        );

    \I__12052\ : LocalMux
    port map (
            O => \N__52459\,
            I => \N__52451\
        );

    \I__12051\ : LocalMux
    port map (
            O => \N__52456\,
            I => \N__52448\
        );

    \I__12050\ : InMux
    port map (
            O => \N__52455\,
            I => \N__52445\
        );

    \I__12049\ : InMux
    port map (
            O => \N__52454\,
            I => \N__52442\
        );

    \I__12048\ : Span4Mux_v
    port map (
            O => \N__52451\,
            I => \N__52439\
        );

    \I__12047\ : Span4Mux_v
    port map (
            O => \N__52448\,
            I => \N__52432\
        );

    \I__12046\ : LocalMux
    port map (
            O => \N__52445\,
            I => \N__52432\
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__52442\,
            I => \N__52432\
        );

    \I__12044\ : Odrv4
    port map (
            O => \N__52439\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__12043\ : Odrv4
    port map (
            O => \N__52432\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__12042\ : InMux
    port map (
            O => \N__52427\,
            I => \N__52413\
        );

    \I__12041\ : InMux
    port map (
            O => \N__52426\,
            I => \N__52408\
        );

    \I__12040\ : InMux
    port map (
            O => \N__52425\,
            I => \N__52408\
        );

    \I__12039\ : InMux
    port map (
            O => \N__52424\,
            I => \N__52405\
        );

    \I__12038\ : InMux
    port map (
            O => \N__52423\,
            I => \N__52402\
        );

    \I__12037\ : InMux
    port map (
            O => \N__52422\,
            I => \N__52397\
        );

    \I__12036\ : InMux
    port map (
            O => \N__52421\,
            I => \N__52394\
        );

    \I__12035\ : InMux
    port map (
            O => \N__52420\,
            I => \N__52389\
        );

    \I__12034\ : InMux
    port map (
            O => \N__52419\,
            I => \N__52389\
        );

    \I__12033\ : CascadeMux
    port map (
            O => \N__52418\,
            I => \N__52384\
        );

    \I__12032\ : InMux
    port map (
            O => \N__52417\,
            I => \N__52379\
        );

    \I__12031\ : InMux
    port map (
            O => \N__52416\,
            I => \N__52379\
        );

    \I__12030\ : LocalMux
    port map (
            O => \N__52413\,
            I => \N__52376\
        );

    \I__12029\ : LocalMux
    port map (
            O => \N__52408\,
            I => \N__52358\
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__52405\,
            I => \N__52355\
        );

    \I__12027\ : LocalMux
    port map (
            O => \N__52402\,
            I => \N__52352\
        );

    \I__12026\ : InMux
    port map (
            O => \N__52401\,
            I => \N__52347\
        );

    \I__12025\ : InMux
    port map (
            O => \N__52400\,
            I => \N__52347\
        );

    \I__12024\ : LocalMux
    port map (
            O => \N__52397\,
            I => \N__52344\
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__52394\,
            I => \N__52339\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__52389\,
            I => \N__52339\
        );

    \I__12021\ : InMux
    port map (
            O => \N__52388\,
            I => \N__52332\
        );

    \I__12020\ : InMux
    port map (
            O => \N__52387\,
            I => \N__52332\
        );

    \I__12019\ : InMux
    port map (
            O => \N__52384\,
            I => \N__52332\
        );

    \I__12018\ : LocalMux
    port map (
            O => \N__52379\,
            I => \N__52329\
        );

    \I__12017\ : Span4Mux_v
    port map (
            O => \N__52376\,
            I => \N__52326\
        );

    \I__12016\ : InMux
    port map (
            O => \N__52375\,
            I => \N__52323\
        );

    \I__12015\ : InMux
    port map (
            O => \N__52374\,
            I => \N__52320\
        );

    \I__12014\ : InMux
    port map (
            O => \N__52373\,
            I => \N__52307\
        );

    \I__12013\ : InMux
    port map (
            O => \N__52372\,
            I => \N__52307\
        );

    \I__12012\ : InMux
    port map (
            O => \N__52371\,
            I => \N__52307\
        );

    \I__12011\ : InMux
    port map (
            O => \N__52370\,
            I => \N__52307\
        );

    \I__12010\ : InMux
    port map (
            O => \N__52369\,
            I => \N__52307\
        );

    \I__12009\ : InMux
    port map (
            O => \N__52368\,
            I => \N__52307\
        );

    \I__12008\ : InMux
    port map (
            O => \N__52367\,
            I => \N__52304\
        );

    \I__12007\ : InMux
    port map (
            O => \N__52366\,
            I => \N__52291\
        );

    \I__12006\ : InMux
    port map (
            O => \N__52365\,
            I => \N__52291\
        );

    \I__12005\ : InMux
    port map (
            O => \N__52364\,
            I => \N__52291\
        );

    \I__12004\ : InMux
    port map (
            O => \N__52363\,
            I => \N__52291\
        );

    \I__12003\ : InMux
    port map (
            O => \N__52362\,
            I => \N__52291\
        );

    \I__12002\ : InMux
    port map (
            O => \N__52361\,
            I => \N__52291\
        );

    \I__12001\ : Span4Mux_h
    port map (
            O => \N__52358\,
            I => \N__52284\
        );

    \I__12000\ : Span4Mux_h
    port map (
            O => \N__52355\,
            I => \N__52284\
        );

    \I__11999\ : Span4Mux_h
    port map (
            O => \N__52352\,
            I => \N__52284\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__52347\,
            I => \N__52275\
        );

    \I__11997\ : Span4Mux_h
    port map (
            O => \N__52344\,
            I => \N__52275\
        );

    \I__11996\ : Span4Mux_v
    port map (
            O => \N__52339\,
            I => \N__52275\
        );

    \I__11995\ : LocalMux
    port map (
            O => \N__52332\,
            I => \N__52275\
        );

    \I__11994\ : Span4Mux_h
    port map (
            O => \N__52329\,
            I => \N__52268\
        );

    \I__11993\ : Span4Mux_h
    port map (
            O => \N__52326\,
            I => \N__52268\
        );

    \I__11992\ : LocalMux
    port map (
            O => \N__52323\,
            I => \N__52268\
        );

    \I__11991\ : LocalMux
    port map (
            O => \N__52320\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__11990\ : LocalMux
    port map (
            O => \N__52307\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__11989\ : LocalMux
    port map (
            O => \N__52304\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__11988\ : LocalMux
    port map (
            O => \N__52291\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__11987\ : Odrv4
    port map (
            O => \N__52284\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__11986\ : Odrv4
    port map (
            O => \N__52275\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__11985\ : Odrv4
    port map (
            O => \N__52268\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__11984\ : InMux
    port map (
            O => \N__52253\,
            I => \N__52250\
        );

    \I__11983\ : LocalMux
    port map (
            O => \N__52250\,
            I => \N__52247\
        );

    \I__11982\ : Span4Mux_h
    port map (
            O => \N__52247\,
            I => \N__52244\
        );

    \I__11981\ : Odrv4
    port map (
            O => \N__52244\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__11980\ : InMux
    port map (
            O => \N__52241\,
            I => \N__52230\
        );

    \I__11979\ : InMux
    port map (
            O => \N__52240\,
            I => \N__52227\
        );

    \I__11978\ : InMux
    port map (
            O => \N__52239\,
            I => \N__52224\
        );

    \I__11977\ : InMux
    port map (
            O => \N__52238\,
            I => \N__52216\
        );

    \I__11976\ : InMux
    port map (
            O => \N__52237\,
            I => \N__52216\
        );

    \I__11975\ : InMux
    port map (
            O => \N__52236\,
            I => \N__52201\
        );

    \I__11974\ : InMux
    port map (
            O => \N__52235\,
            I => \N__52198\
        );

    \I__11973\ : InMux
    port map (
            O => \N__52234\,
            I => \N__52191\
        );

    \I__11972\ : InMux
    port map (
            O => \N__52233\,
            I => \N__52191\
        );

    \I__11971\ : LocalMux
    port map (
            O => \N__52230\,
            I => \N__52184\
        );

    \I__11970\ : LocalMux
    port map (
            O => \N__52227\,
            I => \N__52181\
        );

    \I__11969\ : LocalMux
    port map (
            O => \N__52224\,
            I => \N__52178\
        );

    \I__11968\ : InMux
    port map (
            O => \N__52223\,
            I => \N__52173\
        );

    \I__11967\ : InMux
    port map (
            O => \N__52222\,
            I => \N__52173\
        );

    \I__11966\ : CEMux
    port map (
            O => \N__52221\,
            I => \N__52170\
        );

    \I__11965\ : LocalMux
    port map (
            O => \N__52216\,
            I => \N__52167\
        );

    \I__11964\ : InMux
    port map (
            O => \N__52215\,
            I => \N__52154\
        );

    \I__11963\ : InMux
    port map (
            O => \N__52214\,
            I => \N__52154\
        );

    \I__11962\ : InMux
    port map (
            O => \N__52213\,
            I => \N__52154\
        );

    \I__11961\ : InMux
    port map (
            O => \N__52212\,
            I => \N__52154\
        );

    \I__11960\ : InMux
    port map (
            O => \N__52211\,
            I => \N__52154\
        );

    \I__11959\ : InMux
    port map (
            O => \N__52210\,
            I => \N__52154\
        );

    \I__11958\ : InMux
    port map (
            O => \N__52209\,
            I => \N__52141\
        );

    \I__11957\ : InMux
    port map (
            O => \N__52208\,
            I => \N__52141\
        );

    \I__11956\ : InMux
    port map (
            O => \N__52207\,
            I => \N__52141\
        );

    \I__11955\ : InMux
    port map (
            O => \N__52206\,
            I => \N__52141\
        );

    \I__11954\ : InMux
    port map (
            O => \N__52205\,
            I => \N__52141\
        );

    \I__11953\ : InMux
    port map (
            O => \N__52204\,
            I => \N__52141\
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__52201\,
            I => \N__52136\
        );

    \I__11951\ : LocalMux
    port map (
            O => \N__52198\,
            I => \N__52136\
        );

    \I__11950\ : InMux
    port map (
            O => \N__52197\,
            I => \N__52131\
        );

    \I__11949\ : InMux
    port map (
            O => \N__52196\,
            I => \N__52131\
        );

    \I__11948\ : LocalMux
    port map (
            O => \N__52191\,
            I => \N__52128\
        );

    \I__11947\ : InMux
    port map (
            O => \N__52190\,
            I => \N__52125\
        );

    \I__11946\ : InMux
    port map (
            O => \N__52189\,
            I => \N__52122\
        );

    \I__11945\ : InMux
    port map (
            O => \N__52188\,
            I => \N__52117\
        );

    \I__11944\ : InMux
    port map (
            O => \N__52187\,
            I => \N__52117\
        );

    \I__11943\ : Span4Mux_h
    port map (
            O => \N__52184\,
            I => \N__52112\
        );

    \I__11942\ : Span4Mux_h
    port map (
            O => \N__52181\,
            I => \N__52112\
        );

    \I__11941\ : Span4Mux_v
    port map (
            O => \N__52178\,
            I => \N__52109\
        );

    \I__11940\ : LocalMux
    port map (
            O => \N__52173\,
            I => \N__52106\
        );

    \I__11939\ : LocalMux
    port map (
            O => \N__52170\,
            I => \N__52095\
        );

    \I__11938\ : Span4Mux_v
    port map (
            O => \N__52167\,
            I => \N__52095\
        );

    \I__11937\ : LocalMux
    port map (
            O => \N__52154\,
            I => \N__52095\
        );

    \I__11936\ : LocalMux
    port map (
            O => \N__52141\,
            I => \N__52095\
        );

    \I__11935\ : Span4Mux_v
    port map (
            O => \N__52136\,
            I => \N__52095\
        );

    \I__11934\ : LocalMux
    port map (
            O => \N__52131\,
            I => \N__52090\
        );

    \I__11933\ : Span12Mux_v
    port map (
            O => \N__52128\,
            I => \N__52090\
        );

    \I__11932\ : LocalMux
    port map (
            O => \N__52125\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__11931\ : LocalMux
    port map (
            O => \N__52122\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__11930\ : LocalMux
    port map (
            O => \N__52117\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__11929\ : Odrv4
    port map (
            O => \N__52112\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__11928\ : Odrv4
    port map (
            O => \N__52109\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__11927\ : Odrv12
    port map (
            O => \N__52106\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__11926\ : Odrv4
    port map (
            O => \N__52095\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__11925\ : Odrv12
    port map (
            O => \N__52090\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__11924\ : CascadeMux
    port map (
            O => \N__52073\,
            I => \N__52069\
        );

    \I__11923\ : CascadeMux
    port map (
            O => \N__52072\,
            I => \N__52065\
        );

    \I__11922\ : InMux
    port map (
            O => \N__52069\,
            I => \N__52062\
        );

    \I__11921\ : InMux
    port map (
            O => \N__52068\,
            I => \N__52059\
        );

    \I__11920\ : InMux
    port map (
            O => \N__52065\,
            I => \N__52055\
        );

    \I__11919\ : LocalMux
    port map (
            O => \N__52062\,
            I => \N__52050\
        );

    \I__11918\ : LocalMux
    port map (
            O => \N__52059\,
            I => \N__52050\
        );

    \I__11917\ : InMux
    port map (
            O => \N__52058\,
            I => \N__52047\
        );

    \I__11916\ : LocalMux
    port map (
            O => \N__52055\,
            I => \N__52044\
        );

    \I__11915\ : Span4Mux_v
    port map (
            O => \N__52050\,
            I => \N__52039\
        );

    \I__11914\ : LocalMux
    port map (
            O => \N__52047\,
            I => \N__52039\
        );

    \I__11913\ : Span4Mux_v
    port map (
            O => \N__52044\,
            I => \N__52036\
        );

    \I__11912\ : Span4Mux_s3_v
    port map (
            O => \N__52039\,
            I => \N__52033\
        );

    \I__11911\ : Span4Mux_h
    port map (
            O => \N__52036\,
            I => \N__52030\
        );

    \I__11910\ : Span4Mux_h
    port map (
            O => \N__52033\,
            I => \N__52027\
        );

    \I__11909\ : Odrv4
    port map (
            O => \N__52030\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__11908\ : Odrv4
    port map (
            O => \N__52027\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__11907\ : InMux
    port map (
            O => \N__52022\,
            I => \N__52016\
        );

    \I__11906\ : InMux
    port map (
            O => \N__52021\,
            I => \N__52016\
        );

    \I__11905\ : LocalMux
    port map (
            O => \N__52016\,
            I => \N__52013\
        );

    \I__11904\ : Odrv4
    port map (
            O => \N__52013\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__11903\ : CascadeMux
    port map (
            O => \N__52010\,
            I => \N__52006\
        );

    \I__11902\ : InMux
    port map (
            O => \N__52009\,
            I => \N__52003\
        );

    \I__11901\ : InMux
    port map (
            O => \N__52006\,
            I => \N__52000\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__52003\,
            I => \N__51995\
        );

    \I__11899\ : LocalMux
    port map (
            O => \N__52000\,
            I => \N__51995\
        );

    \I__11898\ : Span4Mux_h
    port map (
            O => \N__51995\,
            I => \N__51992\
        );

    \I__11897\ : Odrv4
    port map (
            O => \N__51992\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__11896\ : CascadeMux
    port map (
            O => \N__51989\,
            I => \N__51986\
        );

    \I__11895\ : InMux
    port map (
            O => \N__51986\,
            I => \N__51980\
        );

    \I__11894\ : InMux
    port map (
            O => \N__51985\,
            I => \N__51980\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__51980\,
            I => \N__51977\
        );

    \I__11892\ : Odrv12
    port map (
            O => \N__51977\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__11891\ : InMux
    port map (
            O => \N__51974\,
            I => \N__51968\
        );

    \I__11890\ : InMux
    port map (
            O => \N__51973\,
            I => \N__51968\
        );

    \I__11889\ : LocalMux
    port map (
            O => \N__51968\,
            I => \N__51965\
        );

    \I__11888\ : Odrv4
    port map (
            O => \N__51965\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__11887\ : CascadeMux
    port map (
            O => \N__51962\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\
        );

    \I__11886\ : InMux
    port map (
            O => \N__51959\,
            I => \N__51956\
        );

    \I__11885\ : LocalMux
    port map (
            O => \N__51956\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\
        );

    \I__11884\ : InMux
    port map (
            O => \N__51953\,
            I => \N__51950\
        );

    \I__11883\ : LocalMux
    port map (
            O => \N__51950\,
            I => \N__51946\
        );

    \I__11882\ : InMux
    port map (
            O => \N__51949\,
            I => \N__51943\
        );

    \I__11881\ : Span4Mux_v
    port map (
            O => \N__51946\,
            I => \N__51938\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__51943\,
            I => \N__51938\
        );

    \I__11879\ : Odrv4
    port map (
            O => \N__51938\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__11878\ : CascadeMux
    port map (
            O => \N__51935\,
            I => \N__51932\
        );

    \I__11877\ : InMux
    port map (
            O => \N__51932\,
            I => \N__51929\
        );

    \I__11876\ : LocalMux
    port map (
            O => \N__51929\,
            I => \N__51925\
        );

    \I__11875\ : InMux
    port map (
            O => \N__51928\,
            I => \N__51922\
        );

    \I__11874\ : Span4Mux_h
    port map (
            O => \N__51925\,
            I => \N__51919\
        );

    \I__11873\ : LocalMux
    port map (
            O => \N__51922\,
            I => \N__51916\
        );

    \I__11872\ : Odrv4
    port map (
            O => \N__51919\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__11871\ : Odrv4
    port map (
            O => \N__51916\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__11870\ : CascadeMux
    port map (
            O => \N__51911\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\
        );

    \I__11869\ : InMux
    port map (
            O => \N__51908\,
            I => \N__51902\
        );

    \I__11868\ : InMux
    port map (
            O => \N__51907\,
            I => \N__51902\
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__51902\,
            I => \N__51899\
        );

    \I__11866\ : Odrv4
    port map (
            O => \N__51899\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__11865\ : InMux
    port map (
            O => \N__51896\,
            I => \N__51890\
        );

    \I__11864\ : InMux
    port map (
            O => \N__51895\,
            I => \N__51890\
        );

    \I__11863\ : LocalMux
    port map (
            O => \N__51890\,
            I => \N__51887\
        );

    \I__11862\ : Odrv12
    port map (
            O => \N__51887\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__11861\ : CascadeMux
    port map (
            O => \N__51884\,
            I => \N__51881\
        );

    \I__11860\ : InMux
    port map (
            O => \N__51881\,
            I => \N__51878\
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__51878\,
            I => \N__51874\
        );

    \I__11858\ : InMux
    port map (
            O => \N__51877\,
            I => \N__51871\
        );

    \I__11857\ : Span4Mux_v
    port map (
            O => \N__51874\,
            I => \N__51866\
        );

    \I__11856\ : LocalMux
    port map (
            O => \N__51871\,
            I => \N__51866\
        );

    \I__11855\ : Odrv4
    port map (
            O => \N__51866\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__11854\ : InMux
    port map (
            O => \N__51863\,
            I => \N__51860\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__51860\,
            I => \N__51856\
        );

    \I__11852\ : InMux
    port map (
            O => \N__51859\,
            I => \N__51853\
        );

    \I__11851\ : Span4Mux_v
    port map (
            O => \N__51856\,
            I => \N__51850\
        );

    \I__11850\ : LocalMux
    port map (
            O => \N__51853\,
            I => \N__51847\
        );

    \I__11849\ : Odrv4
    port map (
            O => \N__51850\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__11848\ : Odrv4
    port map (
            O => \N__51847\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__11847\ : InMux
    port map (
            O => \N__51842\,
            I => \N__51836\
        );

    \I__11846\ : InMux
    port map (
            O => \N__51841\,
            I => \N__51836\
        );

    \I__11845\ : LocalMux
    port map (
            O => \N__51836\,
            I => \N__51833\
        );

    \I__11844\ : Odrv4
    port map (
            O => \N__51833\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__11843\ : InMux
    port map (
            O => \N__51830\,
            I => \N__51824\
        );

    \I__11842\ : InMux
    port map (
            O => \N__51829\,
            I => \N__51824\
        );

    \I__11841\ : LocalMux
    port map (
            O => \N__51824\,
            I => \N__51821\
        );

    \I__11840\ : Odrv12
    port map (
            O => \N__51821\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__11839\ : CascadeMux
    port map (
            O => \N__51818\,
            I => \N__51815\
        );

    \I__11838\ : InMux
    port map (
            O => \N__51815\,
            I => \N__51810\
        );

    \I__11837\ : InMux
    port map (
            O => \N__51814\,
            I => \N__51805\
        );

    \I__11836\ : InMux
    port map (
            O => \N__51813\,
            I => \N__51805\
        );

    \I__11835\ : LocalMux
    port map (
            O => \N__51810\,
            I => \N__51801\
        );

    \I__11834\ : LocalMux
    port map (
            O => \N__51805\,
            I => \N__51798\
        );

    \I__11833\ : InMux
    port map (
            O => \N__51804\,
            I => \N__51795\
        );

    \I__11832\ : Span4Mux_h
    port map (
            O => \N__51801\,
            I => \N__51790\
        );

    \I__11831\ : Span4Mux_h
    port map (
            O => \N__51798\,
            I => \N__51790\
        );

    \I__11830\ : LocalMux
    port map (
            O => \N__51795\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__11829\ : Odrv4
    port map (
            O => \N__51790\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__11828\ : CascadeMux
    port map (
            O => \N__51785\,
            I => \N__51782\
        );

    \I__11827\ : InMux
    port map (
            O => \N__51782\,
            I => \N__51777\
        );

    \I__11826\ : InMux
    port map (
            O => \N__51781\,
            I => \N__51772\
        );

    \I__11825\ : InMux
    port map (
            O => \N__51780\,
            I => \N__51772\
        );

    \I__11824\ : LocalMux
    port map (
            O => \N__51777\,
            I => \N__51768\
        );

    \I__11823\ : LocalMux
    port map (
            O => \N__51772\,
            I => \N__51765\
        );

    \I__11822\ : InMux
    port map (
            O => \N__51771\,
            I => \N__51762\
        );

    \I__11821\ : Span4Mux_h
    port map (
            O => \N__51768\,
            I => \N__51757\
        );

    \I__11820\ : Span4Mux_h
    port map (
            O => \N__51765\,
            I => \N__51757\
        );

    \I__11819\ : LocalMux
    port map (
            O => \N__51762\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__11818\ : Odrv4
    port map (
            O => \N__51757\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__11817\ : CascadeMux
    port map (
            O => \N__51752\,
            I => \N__51749\
        );

    \I__11816\ : InMux
    port map (
            O => \N__51749\,
            I => \N__51743\
        );

    \I__11815\ : InMux
    port map (
            O => \N__51748\,
            I => \N__51740\
        );

    \I__11814\ : InMux
    port map (
            O => \N__51747\,
            I => \N__51737\
        );

    \I__11813\ : InMux
    port map (
            O => \N__51746\,
            I => \N__51734\
        );

    \I__11812\ : LocalMux
    port map (
            O => \N__51743\,
            I => \N__51731\
        );

    \I__11811\ : LocalMux
    port map (
            O => \N__51740\,
            I => \N__51728\
        );

    \I__11810\ : LocalMux
    port map (
            O => \N__51737\,
            I => \N__51723\
        );

    \I__11809\ : LocalMux
    port map (
            O => \N__51734\,
            I => \N__51723\
        );

    \I__11808\ : Span4Mux_v
    port map (
            O => \N__51731\,
            I => \N__51720\
        );

    \I__11807\ : Span4Mux_v
    port map (
            O => \N__51728\,
            I => \N__51717\
        );

    \I__11806\ : Span4Mux_h
    port map (
            O => \N__51723\,
            I => \N__51714\
        );

    \I__11805\ : Odrv4
    port map (
            O => \N__51720\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__11804\ : Odrv4
    port map (
            O => \N__51717\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__11803\ : Odrv4
    port map (
            O => \N__51714\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__11802\ : CascadeMux
    port map (
            O => \N__51707\,
            I => \N__51702\
        );

    \I__11801\ : CascadeMux
    port map (
            O => \N__51706\,
            I => \N__51699\
        );

    \I__11800\ : InMux
    port map (
            O => \N__51705\,
            I => \N__51696\
        );

    \I__11799\ : InMux
    port map (
            O => \N__51702\,
            I => \N__51693\
        );

    \I__11798\ : InMux
    port map (
            O => \N__51699\,
            I => \N__51690\
        );

    \I__11797\ : LocalMux
    port map (
            O => \N__51696\,
            I => \N__51684\
        );

    \I__11796\ : LocalMux
    port map (
            O => \N__51693\,
            I => \N__51684\
        );

    \I__11795\ : LocalMux
    port map (
            O => \N__51690\,
            I => \N__51681\
        );

    \I__11794\ : InMux
    port map (
            O => \N__51689\,
            I => \N__51678\
        );

    \I__11793\ : Span4Mux_h
    port map (
            O => \N__51684\,
            I => \N__51675\
        );

    \I__11792\ : Odrv4
    port map (
            O => \N__51681\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__11791\ : LocalMux
    port map (
            O => \N__51678\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__11790\ : Odrv4
    port map (
            O => \N__51675\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__11789\ : CascadeMux
    port map (
            O => \N__51668\,
            I => \N__51665\
        );

    \I__11788\ : InMux
    port map (
            O => \N__51665\,
            I => \N__51661\
        );

    \I__11787\ : InMux
    port map (
            O => \N__51664\,
            I => \N__51657\
        );

    \I__11786\ : LocalMux
    port map (
            O => \N__51661\,
            I => \N__51653\
        );

    \I__11785\ : InMux
    port map (
            O => \N__51660\,
            I => \N__51650\
        );

    \I__11784\ : LocalMux
    port map (
            O => \N__51657\,
            I => \N__51647\
        );

    \I__11783\ : InMux
    port map (
            O => \N__51656\,
            I => \N__51644\
        );

    \I__11782\ : Span4Mux_h
    port map (
            O => \N__51653\,
            I => \N__51641\
        );

    \I__11781\ : LocalMux
    port map (
            O => \N__51650\,
            I => \N__51638\
        );

    \I__11780\ : Odrv12
    port map (
            O => \N__51647\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__11779\ : LocalMux
    port map (
            O => \N__51644\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__11778\ : Odrv4
    port map (
            O => \N__51641\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__11777\ : Odrv4
    port map (
            O => \N__51638\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__11776\ : InMux
    port map (
            O => \N__51629\,
            I => \N__51623\
        );

    \I__11775\ : InMux
    port map (
            O => \N__51628\,
            I => \N__51623\
        );

    \I__11774\ : LocalMux
    port map (
            O => \N__51623\,
            I => \N__51619\
        );

    \I__11773\ : InMux
    port map (
            O => \N__51622\,
            I => \N__51615\
        );

    \I__11772\ : Span4Mux_v
    port map (
            O => \N__51619\,
            I => \N__51612\
        );

    \I__11771\ : InMux
    port map (
            O => \N__51618\,
            I => \N__51609\
        );

    \I__11770\ : LocalMux
    port map (
            O => \N__51615\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__11769\ : Odrv4
    port map (
            O => \N__51612\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__11768\ : LocalMux
    port map (
            O => \N__51609\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__11767\ : CascadeMux
    port map (
            O => \N__51602\,
            I => \N__51599\
        );

    \I__11766\ : InMux
    port map (
            O => \N__51599\,
            I => \N__51596\
        );

    \I__11765\ : LocalMux
    port map (
            O => \N__51596\,
            I => \N__51590\
        );

    \I__11764\ : InMux
    port map (
            O => \N__51595\,
            I => \N__51587\
        );

    \I__11763\ : InMux
    port map (
            O => \N__51594\,
            I => \N__51582\
        );

    \I__11762\ : InMux
    port map (
            O => \N__51593\,
            I => \N__51582\
        );

    \I__11761\ : Span4Mux_v
    port map (
            O => \N__51590\,
            I => \N__51579\
        );

    \I__11760\ : LocalMux
    port map (
            O => \N__51587\,
            I => \N__51576\
        );

    \I__11759\ : LocalMux
    port map (
            O => \N__51582\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__11758\ : Odrv4
    port map (
            O => \N__51579\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__11757\ : Odrv12
    port map (
            O => \N__51576\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__11756\ : CascadeMux
    port map (
            O => \N__51569\,
            I => \N__51566\
        );

    \I__11755\ : InMux
    port map (
            O => \N__51566\,
            I => \N__51563\
        );

    \I__11754\ : LocalMux
    port map (
            O => \N__51563\,
            I => \N__51559\
        );

    \I__11753\ : CascadeMux
    port map (
            O => \N__51562\,
            I => \N__51556\
        );

    \I__11752\ : Span4Mux_v
    port map (
            O => \N__51559\,
            I => \N__51552\
        );

    \I__11751\ : InMux
    port map (
            O => \N__51556\,
            I => \N__51549\
        );

    \I__11750\ : InMux
    port map (
            O => \N__51555\,
            I => \N__51546\
        );

    \I__11749\ : Odrv4
    port map (
            O => \N__51552\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__51549\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__51546\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__11746\ : InMux
    port map (
            O => \N__51539\,
            I => \N__51536\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__51536\,
            I => \N__51531\
        );

    \I__11744\ : CascadeMux
    port map (
            O => \N__51535\,
            I => \N__51528\
        );

    \I__11743\ : InMux
    port map (
            O => \N__51534\,
            I => \N__51525\
        );

    \I__11742\ : Span4Mux_h
    port map (
            O => \N__51531\,
            I => \N__51522\
        );

    \I__11741\ : InMux
    port map (
            O => \N__51528\,
            I => \N__51519\
        );

    \I__11740\ : LocalMux
    port map (
            O => \N__51525\,
            I => \N__51515\
        );

    \I__11739\ : Span4Mux_v
    port map (
            O => \N__51522\,
            I => \N__51510\
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__51519\,
            I => \N__51510\
        );

    \I__11737\ : InMux
    port map (
            O => \N__51518\,
            I => \N__51507\
        );

    \I__11736\ : Odrv4
    port map (
            O => \N__51515\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__11735\ : Odrv4
    port map (
            O => \N__51510\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__11734\ : LocalMux
    port map (
            O => \N__51507\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__11733\ : CascadeMux
    port map (
            O => \N__51500\,
            I => \N__51497\
        );

    \I__11732\ : InMux
    port map (
            O => \N__51497\,
            I => \N__51492\
        );

    \I__11731\ : InMux
    port map (
            O => \N__51496\,
            I => \N__51489\
        );

    \I__11730\ : InMux
    port map (
            O => \N__51495\,
            I => \N__51486\
        );

    \I__11729\ : LocalMux
    port map (
            O => \N__51492\,
            I => \N__51483\
        );

    \I__11728\ : LocalMux
    port map (
            O => \N__51489\,
            I => \N__51478\
        );

    \I__11727\ : LocalMux
    port map (
            O => \N__51486\,
            I => \N__51478\
        );

    \I__11726\ : Span4Mux_h
    port map (
            O => \N__51483\,
            I => \N__51475\
        );

    \I__11725\ : Span12Mux_s8_v
    port map (
            O => \N__51478\,
            I => \N__51471\
        );

    \I__11724\ : Span4Mux_h
    port map (
            O => \N__51475\,
            I => \N__51468\
        );

    \I__11723\ : InMux
    port map (
            O => \N__51474\,
            I => \N__51465\
        );

    \I__11722\ : Odrv12
    port map (
            O => \N__51471\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__11721\ : Odrv4
    port map (
            O => \N__51468\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__11720\ : LocalMux
    port map (
            O => \N__51465\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__11719\ : CascadeMux
    port map (
            O => \N__51458\,
            I => \current_shift_inst.PI_CTRL.N_77_cascade_\
        );

    \I__11718\ : InMux
    port map (
            O => \N__51455\,
            I => \N__51452\
        );

    \I__11717\ : LocalMux
    port map (
            O => \N__51452\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\
        );

    \I__11716\ : InMux
    port map (
            O => \N__51449\,
            I => \N__51446\
        );

    \I__11715\ : LocalMux
    port map (
            O => \N__51446\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__11714\ : CascadeMux
    port map (
            O => \N__51443\,
            I => \N__51440\
        );

    \I__11713\ : InMux
    port map (
            O => \N__51440\,
            I => \N__51437\
        );

    \I__11712\ : LocalMux
    port map (
            O => \N__51437\,
            I => \N__51433\
        );

    \I__11711\ : InMux
    port map (
            O => \N__51436\,
            I => \N__51428\
        );

    \I__11710\ : Span4Mux_h
    port map (
            O => \N__51433\,
            I => \N__51425\
        );

    \I__11709\ : InMux
    port map (
            O => \N__51432\,
            I => \N__51422\
        );

    \I__11708\ : InMux
    port map (
            O => \N__51431\,
            I => \N__51419\
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__51428\,
            I => \N__51416\
        );

    \I__11706\ : Odrv4
    port map (
            O => \N__51425\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__51422\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__51419\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__11703\ : Odrv12
    port map (
            O => \N__51416\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__11702\ : InMux
    port map (
            O => \N__51407\,
            I => \N__51404\
        );

    \I__11701\ : LocalMux
    port map (
            O => \N__51404\,
            I => \current_shift_inst.PI_CTRL.N_46_16\
        );

    \I__11700\ : InMux
    port map (
            O => \N__51401\,
            I => \N__51398\
        );

    \I__11699\ : LocalMux
    port map (
            O => \N__51398\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\
        );

    \I__11698\ : InMux
    port map (
            O => \N__51395\,
            I => \N__51392\
        );

    \I__11697\ : LocalMux
    port map (
            O => \N__51392\,
            I => \N__51389\
        );

    \I__11696\ : Span4Mux_s3_v
    port map (
            O => \N__51389\,
            I => \N__51386\
        );

    \I__11695\ : Odrv4
    port map (
            O => \N__51386\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__11694\ : CascadeMux
    port map (
            O => \N__51383\,
            I => \N__51380\
        );

    \I__11693\ : InMux
    port map (
            O => \N__51380\,
            I => \N__51374\
        );

    \I__11692\ : InMux
    port map (
            O => \N__51379\,
            I => \N__51371\
        );

    \I__11691\ : InMux
    port map (
            O => \N__51378\,
            I => \N__51368\
        );

    \I__11690\ : CascadeMux
    port map (
            O => \N__51377\,
            I => \N__51365\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__51374\,
            I => \N__51362\
        );

    \I__11688\ : LocalMux
    port map (
            O => \N__51371\,
            I => \N__51359\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__51368\,
            I => \N__51356\
        );

    \I__11686\ : InMux
    port map (
            O => \N__51365\,
            I => \N__51353\
        );

    \I__11685\ : Span4Mux_v
    port map (
            O => \N__51362\,
            I => \N__51346\
        );

    \I__11684\ : Span4Mux_h
    port map (
            O => \N__51359\,
            I => \N__51346\
        );

    \I__11683\ : Span4Mux_v
    port map (
            O => \N__51356\,
            I => \N__51346\
        );

    \I__11682\ : LocalMux
    port map (
            O => \N__51353\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__11681\ : Odrv4
    port map (
            O => \N__51346\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__11680\ : InMux
    port map (
            O => \N__51341\,
            I => \N__51338\
        );

    \I__11679\ : LocalMux
    port map (
            O => \N__51338\,
            I => \N__51335\
        );

    \I__11678\ : Odrv12
    port map (
            O => \N__51335\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__11677\ : CascadeMux
    port map (
            O => \N__51332\,
            I => \N__51328\
        );

    \I__11676\ : CascadeMux
    port map (
            O => \N__51331\,
            I => \N__51325\
        );

    \I__11675\ : InMux
    port map (
            O => \N__51328\,
            I => \N__51321\
        );

    \I__11674\ : InMux
    port map (
            O => \N__51325\,
            I => \N__51316\
        );

    \I__11673\ : InMux
    port map (
            O => \N__51324\,
            I => \N__51316\
        );

    \I__11672\ : LocalMux
    port map (
            O => \N__51321\,
            I => \N__51312\
        );

    \I__11671\ : LocalMux
    port map (
            O => \N__51316\,
            I => \N__51309\
        );

    \I__11670\ : InMux
    port map (
            O => \N__51315\,
            I => \N__51306\
        );

    \I__11669\ : Span4Mux_h
    port map (
            O => \N__51312\,
            I => \N__51301\
        );

    \I__11668\ : Span4Mux_v
    port map (
            O => \N__51309\,
            I => \N__51301\
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__51306\,
            I => \N__51298\
        );

    \I__11666\ : Odrv4
    port map (
            O => \N__51301\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__11665\ : Odrv4
    port map (
            O => \N__51298\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__11664\ : InMux
    port map (
            O => \N__51293\,
            I => \N__51290\
        );

    \I__11663\ : LocalMux
    port map (
            O => \N__51290\,
            I => \N__51287\
        );

    \I__11662\ : Span4Mux_v
    port map (
            O => \N__51287\,
            I => \N__51284\
        );

    \I__11661\ : Odrv4
    port map (
            O => \N__51284\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__11660\ : CascadeMux
    port map (
            O => \N__51281\,
            I => \N__51277\
        );

    \I__11659\ : CascadeMux
    port map (
            O => \N__51280\,
            I => \N__51272\
        );

    \I__11658\ : InMux
    port map (
            O => \N__51277\,
            I => \N__51269\
        );

    \I__11657\ : InMux
    port map (
            O => \N__51276\,
            I => \N__51264\
        );

    \I__11656\ : InMux
    port map (
            O => \N__51275\,
            I => \N__51264\
        );

    \I__11655\ : InMux
    port map (
            O => \N__51272\,
            I => \N__51261\
        );

    \I__11654\ : LocalMux
    port map (
            O => \N__51269\,
            I => \N__51254\
        );

    \I__11653\ : LocalMux
    port map (
            O => \N__51264\,
            I => \N__51254\
        );

    \I__11652\ : LocalMux
    port map (
            O => \N__51261\,
            I => \N__51254\
        );

    \I__11651\ : Span4Mux_v
    port map (
            O => \N__51254\,
            I => \N__51251\
        );

    \I__11650\ : Odrv4
    port map (
            O => \N__51251\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__11649\ : InMux
    port map (
            O => \N__51248\,
            I => \N__51245\
        );

    \I__11648\ : LocalMux
    port map (
            O => \N__51245\,
            I => \N__51242\
        );

    \I__11647\ : Odrv4
    port map (
            O => \N__51242\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\
        );

    \I__11646\ : CascadeMux
    port map (
            O => \N__51239\,
            I => \N__51236\
        );

    \I__11645\ : InMux
    port map (
            O => \N__51236\,
            I => \N__51233\
        );

    \I__11644\ : LocalMux
    port map (
            O => \N__51233\,
            I => \N__51227\
        );

    \I__11643\ : InMux
    port map (
            O => \N__51232\,
            I => \N__51224\
        );

    \I__11642\ : InMux
    port map (
            O => \N__51231\,
            I => \N__51219\
        );

    \I__11641\ : InMux
    port map (
            O => \N__51230\,
            I => \N__51219\
        );

    \I__11640\ : Odrv4
    port map (
            O => \N__51227\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__51224\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__11638\ : LocalMux
    port map (
            O => \N__51219\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__11637\ : InMux
    port map (
            O => \N__51212\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__11636\ : InMux
    port map (
            O => \N__51209\,
            I => \N__51206\
        );

    \I__11635\ : LocalMux
    port map (
            O => \N__51206\,
            I => \N__51203\
        );

    \I__11634\ : Odrv4
    port map (
            O => \N__51203\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\
        );

    \I__11633\ : CascadeMux
    port map (
            O => \N__51200\,
            I => \N__51197\
        );

    \I__11632\ : InMux
    port map (
            O => \N__51197\,
            I => \N__51193\
        );

    \I__11631\ : CascadeMux
    port map (
            O => \N__51196\,
            I => \N__51190\
        );

    \I__11630\ : LocalMux
    port map (
            O => \N__51193\,
            I => \N__51185\
        );

    \I__11629\ : InMux
    port map (
            O => \N__51190\,
            I => \N__51182\
        );

    \I__11628\ : InMux
    port map (
            O => \N__51189\,
            I => \N__51179\
        );

    \I__11627\ : InMux
    port map (
            O => \N__51188\,
            I => \N__51176\
        );

    \I__11626\ : Odrv4
    port map (
            O => \N__51185\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__51182\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__11624\ : LocalMux
    port map (
            O => \N__51179\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__11623\ : LocalMux
    port map (
            O => \N__51176\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__11622\ : InMux
    port map (
            O => \N__51167\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__11621\ : InMux
    port map (
            O => \N__51164\,
            I => \N__51161\
        );

    \I__11620\ : LocalMux
    port map (
            O => \N__51161\,
            I => \N__51158\
        );

    \I__11619\ : Span4Mux_v
    port map (
            O => \N__51158\,
            I => \N__51155\
        );

    \I__11618\ : Odrv4
    port map (
            O => \N__51155\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\
        );

    \I__11617\ : CascadeMux
    port map (
            O => \N__51152\,
            I => \N__51149\
        );

    \I__11616\ : InMux
    port map (
            O => \N__51149\,
            I => \N__51145\
        );

    \I__11615\ : CascadeMux
    port map (
            O => \N__51148\,
            I => \N__51142\
        );

    \I__11614\ : LocalMux
    port map (
            O => \N__51145\,
            I => \N__51137\
        );

    \I__11613\ : InMux
    port map (
            O => \N__51142\,
            I => \N__51134\
        );

    \I__11612\ : InMux
    port map (
            O => \N__51141\,
            I => \N__51131\
        );

    \I__11611\ : InMux
    port map (
            O => \N__51140\,
            I => \N__51128\
        );

    \I__11610\ : Odrv12
    port map (
            O => \N__51137\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__11609\ : LocalMux
    port map (
            O => \N__51134\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__11608\ : LocalMux
    port map (
            O => \N__51131\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__11607\ : LocalMux
    port map (
            O => \N__51128\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__11606\ : InMux
    port map (
            O => \N__51119\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__11605\ : InMux
    port map (
            O => \N__51116\,
            I => \N__51113\
        );

    \I__11604\ : LocalMux
    port map (
            O => \N__51113\,
            I => \N__51110\
        );

    \I__11603\ : Span4Mux_h
    port map (
            O => \N__51110\,
            I => \N__51107\
        );

    \I__11602\ : Odrv4
    port map (
            O => \N__51107\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\
        );

    \I__11601\ : CascadeMux
    port map (
            O => \N__51104\,
            I => \N__51101\
        );

    \I__11600\ : InMux
    port map (
            O => \N__51101\,
            I => \N__51097\
        );

    \I__11599\ : CascadeMux
    port map (
            O => \N__51100\,
            I => \N__51093\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__51097\,
            I => \N__51089\
        );

    \I__11597\ : InMux
    port map (
            O => \N__51096\,
            I => \N__51086\
        );

    \I__11596\ : InMux
    port map (
            O => \N__51093\,
            I => \N__51081\
        );

    \I__11595\ : InMux
    port map (
            O => \N__51092\,
            I => \N__51081\
        );

    \I__11594\ : Odrv12
    port map (
            O => \N__51089\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__51086\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__11592\ : LocalMux
    port map (
            O => \N__51081\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__11591\ : InMux
    port map (
            O => \N__51074\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__11590\ : InMux
    port map (
            O => \N__51071\,
            I => \N__51067\
        );

    \I__11589\ : CascadeMux
    port map (
            O => \N__51070\,
            I => \N__51064\
        );

    \I__11588\ : LocalMux
    port map (
            O => \N__51067\,
            I => \N__51059\
        );

    \I__11587\ : InMux
    port map (
            O => \N__51064\,
            I => \N__51056\
        );

    \I__11586\ : InMux
    port map (
            O => \N__51063\,
            I => \N__51053\
        );

    \I__11585\ : InMux
    port map (
            O => \N__51062\,
            I => \N__51050\
        );

    \I__11584\ : Odrv12
    port map (
            O => \N__51059\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__11583\ : LocalMux
    port map (
            O => \N__51056\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__11582\ : LocalMux
    port map (
            O => \N__51053\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__11581\ : LocalMux
    port map (
            O => \N__51050\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__11580\ : CascadeMux
    port map (
            O => \N__51041\,
            I => \N__51038\
        );

    \I__11579\ : InMux
    port map (
            O => \N__51038\,
            I => \N__51035\
        );

    \I__11578\ : LocalMux
    port map (
            O => \N__51035\,
            I => \N__51032\
        );

    \I__11577\ : Span4Mux_v
    port map (
            O => \N__51032\,
            I => \N__51029\
        );

    \I__11576\ : Odrv4
    port map (
            O => \N__51029\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\
        );

    \I__11575\ : InMux
    port map (
            O => \N__51026\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__11574\ : InMux
    port map (
            O => \N__51023\,
            I => \N__51020\
        );

    \I__11573\ : LocalMux
    port map (
            O => \N__51020\,
            I => \N__51017\
        );

    \I__11572\ : Odrv4
    port map (
            O => \N__51017\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\
        );

    \I__11571\ : InMux
    port map (
            O => \N__51014\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__11570\ : CascadeMux
    port map (
            O => \N__51011\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__11569\ : InMux
    port map (
            O => \N__51008\,
            I => \N__51005\
        );

    \I__11568\ : LocalMux
    port map (
            O => \N__51005\,
            I => \current_shift_inst.PI_CTRL.N_44\
        );

    \I__11567\ : InMux
    port map (
            O => \N__51002\,
            I => \N__50999\
        );

    \I__11566\ : LocalMux
    port map (
            O => \N__50999\,
            I => \N__50996\
        );

    \I__11565\ : Odrv4
    port map (
            O => \N__50996\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__11564\ : InMux
    port map (
            O => \N__50993\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__11563\ : InMux
    port map (
            O => \N__50990\,
            I => \N__50987\
        );

    \I__11562\ : LocalMux
    port map (
            O => \N__50987\,
            I => \N__50984\
        );

    \I__11561\ : Span12Mux_s7_v
    port map (
            O => \N__50984\,
            I => \N__50981\
        );

    \I__11560\ : Odrv12
    port map (
            O => \N__50981\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__11559\ : InMux
    port map (
            O => \N__50978\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__11558\ : InMux
    port map (
            O => \N__50975\,
            I => \N__50972\
        );

    \I__11557\ : LocalMux
    port map (
            O => \N__50972\,
            I => \N__50969\
        );

    \I__11556\ : Odrv4
    port map (
            O => \N__50969\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__11555\ : InMux
    port map (
            O => \N__50966\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__11554\ : InMux
    port map (
            O => \N__50963\,
            I => \N__50960\
        );

    \I__11553\ : LocalMux
    port map (
            O => \N__50960\,
            I => \N__50957\
        );

    \I__11552\ : Odrv4
    port map (
            O => \N__50957\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__11551\ : CascadeMux
    port map (
            O => \N__50954\,
            I => \N__50951\
        );

    \I__11550\ : InMux
    port map (
            O => \N__50951\,
            I => \N__50946\
        );

    \I__11549\ : InMux
    port map (
            O => \N__50950\,
            I => \N__50940\
        );

    \I__11548\ : InMux
    port map (
            O => \N__50949\,
            I => \N__50940\
        );

    \I__11547\ : LocalMux
    port map (
            O => \N__50946\,
            I => \N__50937\
        );

    \I__11546\ : InMux
    port map (
            O => \N__50945\,
            I => \N__50934\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__50940\,
            I => \N__50931\
        );

    \I__11544\ : Odrv4
    port map (
            O => \N__50937\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__11543\ : LocalMux
    port map (
            O => \N__50934\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__11542\ : Odrv4
    port map (
            O => \N__50931\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__11541\ : InMux
    port map (
            O => \N__50924\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__11540\ : CascadeMux
    port map (
            O => \N__50921\,
            I => \N__50918\
        );

    \I__11539\ : InMux
    port map (
            O => \N__50918\,
            I => \N__50915\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__50915\,
            I => \N__50912\
        );

    \I__11537\ : Odrv4
    port map (
            O => \N__50912\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__11536\ : InMux
    port map (
            O => \N__50909\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__11535\ : InMux
    port map (
            O => \N__50906\,
            I => \N__50900\
        );

    \I__11534\ : InMux
    port map (
            O => \N__50905\,
            I => \N__50897\
        );

    \I__11533\ : InMux
    port map (
            O => \N__50904\,
            I => \N__50892\
        );

    \I__11532\ : InMux
    port map (
            O => \N__50903\,
            I => \N__50892\
        );

    \I__11531\ : LocalMux
    port map (
            O => \N__50900\,
            I => \N__50889\
        );

    \I__11530\ : LocalMux
    port map (
            O => \N__50897\,
            I => \N__50884\
        );

    \I__11529\ : LocalMux
    port map (
            O => \N__50892\,
            I => \N__50884\
        );

    \I__11528\ : Odrv4
    port map (
            O => \N__50889\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__11527\ : Odrv4
    port map (
            O => \N__50884\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__11526\ : CascadeMux
    port map (
            O => \N__50879\,
            I => \N__50876\
        );

    \I__11525\ : InMux
    port map (
            O => \N__50876\,
            I => \N__50873\
        );

    \I__11524\ : LocalMux
    port map (
            O => \N__50873\,
            I => \N__50870\
        );

    \I__11523\ : Span4Mux_h
    port map (
            O => \N__50870\,
            I => \N__50867\
        );

    \I__11522\ : Odrv4
    port map (
            O => \N__50867\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__11521\ : InMux
    port map (
            O => \N__50864\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__11520\ : InMux
    port map (
            O => \N__50861\,
            I => \N__50858\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__50858\,
            I => \N__50855\
        );

    \I__11518\ : Span4Mux_h
    port map (
            O => \N__50855\,
            I => \N__50852\
        );

    \I__11517\ : Odrv4
    port map (
            O => \N__50852\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__11516\ : CascadeMux
    port map (
            O => \N__50849\,
            I => \N__50845\
        );

    \I__11515\ : CascadeMux
    port map (
            O => \N__50848\,
            I => \N__50841\
        );

    \I__11514\ : InMux
    port map (
            O => \N__50845\,
            I => \N__50837\
        );

    \I__11513\ : CascadeMux
    port map (
            O => \N__50844\,
            I => \N__50834\
        );

    \I__11512\ : InMux
    port map (
            O => \N__50841\,
            I => \N__50829\
        );

    \I__11511\ : InMux
    port map (
            O => \N__50840\,
            I => \N__50829\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__50837\,
            I => \N__50826\
        );

    \I__11509\ : InMux
    port map (
            O => \N__50834\,
            I => \N__50823\
        );

    \I__11508\ : LocalMux
    port map (
            O => \N__50829\,
            I => \N__50820\
        );

    \I__11507\ : Odrv12
    port map (
            O => \N__50826\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__11506\ : LocalMux
    port map (
            O => \N__50823\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__11505\ : Odrv4
    port map (
            O => \N__50820\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__11504\ : InMux
    port map (
            O => \N__50813\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\
        );

    \I__11503\ : InMux
    port map (
            O => \N__50810\,
            I => \N__50807\
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__50807\,
            I => \N__50804\
        );

    \I__11501\ : Odrv4
    port map (
            O => \N__50804\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__11500\ : CascadeMux
    port map (
            O => \N__50801\,
            I => \N__50798\
        );

    \I__11499\ : InMux
    port map (
            O => \N__50798\,
            I => \N__50795\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__50795\,
            I => \N__50790\
        );

    \I__11497\ : CascadeMux
    port map (
            O => \N__50794\,
            I => \N__50787\
        );

    \I__11496\ : CascadeMux
    port map (
            O => \N__50793\,
            I => \N__50783\
        );

    \I__11495\ : Span4Mux_h
    port map (
            O => \N__50790\,
            I => \N__50780\
        );

    \I__11494\ : InMux
    port map (
            O => \N__50787\,
            I => \N__50777\
        );

    \I__11493\ : InMux
    port map (
            O => \N__50786\,
            I => \N__50772\
        );

    \I__11492\ : InMux
    port map (
            O => \N__50783\,
            I => \N__50772\
        );

    \I__11491\ : Odrv4
    port map (
            O => \N__50780\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__50777\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__11489\ : LocalMux
    port map (
            O => \N__50772\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__11488\ : InMux
    port map (
            O => \N__50765\,
            I => \bfn_18_26_0_\
        );

    \I__11487\ : InMux
    port map (
            O => \N__50762\,
            I => \N__50759\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__50759\,
            I => \N__50756\
        );

    \I__11485\ : Odrv4
    port map (
            O => \N__50756\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__11484\ : CascadeMux
    port map (
            O => \N__50753\,
            I => \N__50750\
        );

    \I__11483\ : InMux
    port map (
            O => \N__50750\,
            I => \N__50744\
        );

    \I__11482\ : InMux
    port map (
            O => \N__50749\,
            I => \N__50741\
        );

    \I__11481\ : InMux
    port map (
            O => \N__50748\,
            I => \N__50736\
        );

    \I__11480\ : InMux
    port map (
            O => \N__50747\,
            I => \N__50736\
        );

    \I__11479\ : LocalMux
    port map (
            O => \N__50744\,
            I => \N__50731\
        );

    \I__11478\ : LocalMux
    port map (
            O => \N__50741\,
            I => \N__50731\
        );

    \I__11477\ : LocalMux
    port map (
            O => \N__50736\,
            I => \N__50728\
        );

    \I__11476\ : Span4Mux_h
    port map (
            O => \N__50731\,
            I => \N__50725\
        );

    \I__11475\ : Odrv4
    port map (
            O => \N__50728\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__11474\ : Odrv4
    port map (
            O => \N__50725\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__11473\ : InMux
    port map (
            O => \N__50720\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__11472\ : InMux
    port map (
            O => \N__50717\,
            I => \N__50714\
        );

    \I__11471\ : LocalMux
    port map (
            O => \N__50714\,
            I => \N__50711\
        );

    \I__11470\ : Odrv12
    port map (
            O => \N__50711\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__11469\ : InMux
    port map (
            O => \N__50708\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__11468\ : InMux
    port map (
            O => \N__50705\,
            I => \N__50702\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__50702\,
            I => \N__50699\
        );

    \I__11466\ : Odrv12
    port map (
            O => \N__50699\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__11465\ : CascadeMux
    port map (
            O => \N__50696\,
            I => \N__50693\
        );

    \I__11464\ : InMux
    port map (
            O => \N__50693\,
            I => \N__50689\
        );

    \I__11463\ : CascadeMux
    port map (
            O => \N__50692\,
            I => \N__50686\
        );

    \I__11462\ : LocalMux
    port map (
            O => \N__50689\,
            I => \N__50682\
        );

    \I__11461\ : InMux
    port map (
            O => \N__50686\,
            I => \N__50678\
        );

    \I__11460\ : InMux
    port map (
            O => \N__50685\,
            I => \N__50675\
        );

    \I__11459\ : Span4Mux_h
    port map (
            O => \N__50682\,
            I => \N__50672\
        );

    \I__11458\ : CascadeMux
    port map (
            O => \N__50681\,
            I => \N__50669\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__50678\,
            I => \N__50664\
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__50675\,
            I => \N__50664\
        );

    \I__11455\ : Span4Mux_v
    port map (
            O => \N__50672\,
            I => \N__50661\
        );

    \I__11454\ : InMux
    port map (
            O => \N__50669\,
            I => \N__50658\
        );

    \I__11453\ : Span12Mux_v
    port map (
            O => \N__50664\,
            I => \N__50655\
        );

    \I__11452\ : Odrv4
    port map (
            O => \N__50661\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__50658\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__11450\ : Odrv12
    port map (
            O => \N__50655\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__11449\ : InMux
    port map (
            O => \N__50648\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__11448\ : InMux
    port map (
            O => \N__50645\,
            I => \N__50642\
        );

    \I__11447\ : LocalMux
    port map (
            O => \N__50642\,
            I => \N__50639\
        );

    \I__11446\ : Odrv12
    port map (
            O => \N__50639\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__11445\ : CascadeMux
    port map (
            O => \N__50636\,
            I => \N__50633\
        );

    \I__11444\ : InMux
    port map (
            O => \N__50633\,
            I => \N__50630\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__50630\,
            I => \N__50626\
        );

    \I__11442\ : InMux
    port map (
            O => \N__50629\,
            I => \N__50623\
        );

    \I__11441\ : Span4Mux_h
    port map (
            O => \N__50626\,
            I => \N__50619\
        );

    \I__11440\ : LocalMux
    port map (
            O => \N__50623\,
            I => \N__50615\
        );

    \I__11439\ : InMux
    port map (
            O => \N__50622\,
            I => \N__50612\
        );

    \I__11438\ : Span4Mux_v
    port map (
            O => \N__50619\,
            I => \N__50609\
        );

    \I__11437\ : InMux
    port map (
            O => \N__50618\,
            I => \N__50606\
        );

    \I__11436\ : Span4Mux_v
    port map (
            O => \N__50615\,
            I => \N__50603\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__50612\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__11434\ : Odrv4
    port map (
            O => \N__50609\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__50606\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__11432\ : Odrv4
    port map (
            O => \N__50603\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__11431\ : InMux
    port map (
            O => \N__50594\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__11430\ : InMux
    port map (
            O => \N__50591\,
            I => \N__50588\
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__50588\,
            I => \N__50585\
        );

    \I__11428\ : Odrv4
    port map (
            O => \N__50585\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__11427\ : CascadeMux
    port map (
            O => \N__50582\,
            I => \N__50579\
        );

    \I__11426\ : InMux
    port map (
            O => \N__50579\,
            I => \N__50575\
        );

    \I__11425\ : InMux
    port map (
            O => \N__50578\,
            I => \N__50572\
        );

    \I__11424\ : LocalMux
    port map (
            O => \N__50575\,
            I => \N__50565\
        );

    \I__11423\ : LocalMux
    port map (
            O => \N__50572\,
            I => \N__50565\
        );

    \I__11422\ : InMux
    port map (
            O => \N__50571\,
            I => \N__50562\
        );

    \I__11421\ : InMux
    port map (
            O => \N__50570\,
            I => \N__50559\
        );

    \I__11420\ : Span4Mux_h
    port map (
            O => \N__50565\,
            I => \N__50556\
        );

    \I__11419\ : LocalMux
    port map (
            O => \N__50562\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__50559\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__11417\ : Odrv4
    port map (
            O => \N__50556\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__11416\ : InMux
    port map (
            O => \N__50549\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__11415\ : InMux
    port map (
            O => \N__50546\,
            I => \N__50543\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__50543\,
            I => \N__50540\
        );

    \I__11413\ : Span4Mux_h
    port map (
            O => \N__50540\,
            I => \N__50537\
        );

    \I__11412\ : Odrv4
    port map (
            O => \N__50537\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__11411\ : CascadeMux
    port map (
            O => \N__50534\,
            I => \N__50531\
        );

    \I__11410\ : InMux
    port map (
            O => \N__50531\,
            I => \N__50528\
        );

    \I__11409\ : LocalMux
    port map (
            O => \N__50528\,
            I => \N__50523\
        );

    \I__11408\ : InMux
    port map (
            O => \N__50527\,
            I => \N__50517\
        );

    \I__11407\ : InMux
    port map (
            O => \N__50526\,
            I => \N__50517\
        );

    \I__11406\ : Span4Mux_v
    port map (
            O => \N__50523\,
            I => \N__50514\
        );

    \I__11405\ : InMux
    port map (
            O => \N__50522\,
            I => \N__50511\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__50517\,
            I => \N__50508\
        );

    \I__11403\ : Odrv4
    port map (
            O => \N__50514\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__11402\ : LocalMux
    port map (
            O => \N__50511\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__11401\ : Odrv4
    port map (
            O => \N__50508\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__11400\ : InMux
    port map (
            O => \N__50501\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__11399\ : InMux
    port map (
            O => \N__50498\,
            I => \N__50495\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__50495\,
            I => \N__50492\
        );

    \I__11397\ : Odrv12
    port map (
            O => \N__50492\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__11396\ : InMux
    port map (
            O => \N__50489\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\
        );

    \I__11395\ : InMux
    port map (
            O => \N__50486\,
            I => \N__50483\
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__50483\,
            I => \N__50480\
        );

    \I__11393\ : Span4Mux_h
    port map (
            O => \N__50480\,
            I => \N__50477\
        );

    \I__11392\ : Span4Mux_h
    port map (
            O => \N__50477\,
            I => \N__50474\
        );

    \I__11391\ : Odrv4
    port map (
            O => \N__50474\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__11390\ : InMux
    port map (
            O => \N__50471\,
            I => \bfn_18_25_0_\
        );

    \I__11389\ : InMux
    port map (
            O => \N__50468\,
            I => \N__50465\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__50465\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__11387\ : InMux
    port map (
            O => \N__50462\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__11386\ : CascadeMux
    port map (
            O => \N__50459\,
            I => \N__50456\
        );

    \I__11385\ : InMux
    port map (
            O => \N__50456\,
            I => \N__50453\
        );

    \I__11384\ : LocalMux
    port map (
            O => \N__50453\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__11383\ : InMux
    port map (
            O => \N__50450\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__11382\ : InMux
    port map (
            O => \N__50447\,
            I => \N__50444\
        );

    \I__11381\ : LocalMux
    port map (
            O => \N__50444\,
            I => \N__50441\
        );

    \I__11380\ : Odrv4
    port map (
            O => \N__50441\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__11379\ : InMux
    port map (
            O => \N__50438\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__11378\ : InMux
    port map (
            O => \N__50435\,
            I => \N__50432\
        );

    \I__11377\ : LocalMux
    port map (
            O => \N__50432\,
            I => \N__50429\
        );

    \I__11376\ : Span4Mux_h
    port map (
            O => \N__50429\,
            I => \N__50426\
        );

    \I__11375\ : Odrv4
    port map (
            O => \N__50426\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__11374\ : InMux
    port map (
            O => \N__50423\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__11373\ : InMux
    port map (
            O => \N__50420\,
            I => \N__50417\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__50417\,
            I => \N__50414\
        );

    \I__11371\ : Odrv12
    port map (
            O => \N__50414\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__11370\ : InMux
    port map (
            O => \N__50411\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__11369\ : InMux
    port map (
            O => \N__50408\,
            I => \N__50405\
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__50405\,
            I => \N__50402\
        );

    \I__11367\ : Odrv12
    port map (
            O => \N__50402\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__11366\ : InMux
    port map (
            O => \N__50399\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__11365\ : InMux
    port map (
            O => \N__50396\,
            I => \N__50393\
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__50393\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__11363\ : InMux
    port map (
            O => \N__50390\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\
        );

    \I__11362\ : InMux
    port map (
            O => \N__50387\,
            I => \N__50384\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__50384\,
            I => \N__50381\
        );

    \I__11360\ : Odrv4
    port map (
            O => \N__50381\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__11359\ : InMux
    port map (
            O => \N__50378\,
            I => \bfn_18_24_0_\
        );

    \I__11358\ : InMux
    port map (
            O => \N__50375\,
            I => \N__50371\
        );

    \I__11357\ : InMux
    port map (
            O => \N__50374\,
            I => \N__50368\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__50371\,
            I => \N__50365\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__50368\,
            I => \N__50360\
        );

    \I__11354\ : Span12Mux_s8_v
    port map (
            O => \N__50365\,
            I => \N__50360\
        );

    \I__11353\ : Odrv12
    port map (
            O => \N__50360\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__11352\ : InMux
    port map (
            O => \N__50357\,
            I => \N__50354\
        );

    \I__11351\ : LocalMux
    port map (
            O => \N__50354\,
            I => \N__50350\
        );

    \I__11350\ : InMux
    port map (
            O => \N__50353\,
            I => \N__50347\
        );

    \I__11349\ : Span4Mux_v
    port map (
            O => \N__50350\,
            I => \N__50344\
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__50347\,
            I => \N__50339\
        );

    \I__11347\ : Span4Mux_h
    port map (
            O => \N__50344\,
            I => \N__50339\
        );

    \I__11346\ : Span4Mux_h
    port map (
            O => \N__50339\,
            I => \N__50336\
        );

    \I__11345\ : Odrv4
    port map (
            O => \N__50336\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__11344\ : InMux
    port map (
            O => \N__50333\,
            I => \N__50330\
        );

    \I__11343\ : LocalMux
    port map (
            O => \N__50330\,
            I => \N__50326\
        );

    \I__11342\ : InMux
    port map (
            O => \N__50329\,
            I => \N__50323\
        );

    \I__11341\ : Span4Mux_s2_h
    port map (
            O => \N__50326\,
            I => \N__50320\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__50323\,
            I => \N__50315\
        );

    \I__11339\ : Span4Mux_h
    port map (
            O => \N__50320\,
            I => \N__50315\
        );

    \I__11338\ : Span4Mux_v
    port map (
            O => \N__50315\,
            I => \N__50312\
        );

    \I__11337\ : Odrv4
    port map (
            O => \N__50312\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__11336\ : InMux
    port map (
            O => \N__50309\,
            I => \N__50306\
        );

    \I__11335\ : LocalMux
    port map (
            O => \N__50306\,
            I => \N__50303\
        );

    \I__11334\ : Span4Mux_s1_h
    port map (
            O => \N__50303\,
            I => \N__50299\
        );

    \I__11333\ : InMux
    port map (
            O => \N__50302\,
            I => \N__50296\
        );

    \I__11332\ : Span4Mux_h
    port map (
            O => \N__50299\,
            I => \N__50293\
        );

    \I__11331\ : LocalMux
    port map (
            O => \N__50296\,
            I => \N__50290\
        );

    \I__11330\ : Span4Mux_h
    port map (
            O => \N__50293\,
            I => \N__50287\
        );

    \I__11329\ : Odrv4
    port map (
            O => \N__50290\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__11328\ : Odrv4
    port map (
            O => \N__50287\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__11327\ : InMux
    port map (
            O => \N__50282\,
            I => \N__50279\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__50279\,
            I => \N__50275\
        );

    \I__11325\ : InMux
    port map (
            O => \N__50278\,
            I => \N__50272\
        );

    \I__11324\ : Span4Mux_v
    port map (
            O => \N__50275\,
            I => \N__50269\
        );

    \I__11323\ : LocalMux
    port map (
            O => \N__50272\,
            I => \N__50264\
        );

    \I__11322\ : Span4Mux_h
    port map (
            O => \N__50269\,
            I => \N__50264\
        );

    \I__11321\ : Span4Mux_h
    port map (
            O => \N__50264\,
            I => \N__50261\
        );

    \I__11320\ : Odrv4
    port map (
            O => \N__50261\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__11319\ : InMux
    port map (
            O => \N__50258\,
            I => \N__50254\
        );

    \I__11318\ : InMux
    port map (
            O => \N__50257\,
            I => \N__50251\
        );

    \I__11317\ : LocalMux
    port map (
            O => \N__50254\,
            I => \N__50248\
        );

    \I__11316\ : LocalMux
    port map (
            O => \N__50251\,
            I => \N__50245\
        );

    \I__11315\ : Span12Mux_s10_h
    port map (
            O => \N__50248\,
            I => \N__50242\
        );

    \I__11314\ : Odrv4
    port map (
            O => \N__50245\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__11313\ : Odrv12
    port map (
            O => \N__50242\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__11312\ : InMux
    port map (
            O => \N__50237\,
            I => \N__50234\
        );

    \I__11311\ : LocalMux
    port map (
            O => \N__50234\,
            I => \N__50230\
        );

    \I__11310\ : InMux
    port map (
            O => \N__50233\,
            I => \N__50227\
        );

    \I__11309\ : Span4Mux_s2_h
    port map (
            O => \N__50230\,
            I => \N__50224\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__50227\,
            I => \N__50219\
        );

    \I__11307\ : Span4Mux_h
    port map (
            O => \N__50224\,
            I => \N__50219\
        );

    \I__11306\ : Span4Mux_v
    port map (
            O => \N__50219\,
            I => \N__50216\
        );

    \I__11305\ : Odrv4
    port map (
            O => \N__50216\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__11304\ : InMux
    port map (
            O => \N__50213\,
            I => \N__50210\
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__50210\,
            I => \N__50207\
        );

    \I__11302\ : Span4Mux_s2_h
    port map (
            O => \N__50207\,
            I => \N__50203\
        );

    \I__11301\ : InMux
    port map (
            O => \N__50206\,
            I => \N__50200\
        );

    \I__11300\ : Span4Mux_h
    port map (
            O => \N__50203\,
            I => \N__50197\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__50200\,
            I => \N__50194\
        );

    \I__11298\ : Span4Mux_h
    port map (
            O => \N__50197\,
            I => \N__50191\
        );

    \I__11297\ : Odrv4
    port map (
            O => \N__50194\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__11296\ : Odrv4
    port map (
            O => \N__50191\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__11295\ : InMux
    port map (
            O => \N__50186\,
            I => \N__50182\
        );

    \I__11294\ : InMux
    port map (
            O => \N__50185\,
            I => \N__50179\
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__50182\,
            I => \N__50176\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__50179\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__11291\ : Odrv4
    port map (
            O => \N__50176\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__11290\ : InMux
    port map (
            O => \N__50171\,
            I => \N__50168\
        );

    \I__11289\ : LocalMux
    port map (
            O => \N__50168\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\
        );

    \I__11288\ : InMux
    port map (
            O => \N__50165\,
            I => \N__50159\
        );

    \I__11287\ : InMux
    port map (
            O => \N__50164\,
            I => \N__50159\
        );

    \I__11286\ : LocalMux
    port map (
            O => \N__50159\,
            I => \N__50155\
        );

    \I__11285\ : InMux
    port map (
            O => \N__50158\,
            I => \N__50152\
        );

    \I__11284\ : Span4Mux_v
    port map (
            O => \N__50155\,
            I => \N__50149\
        );

    \I__11283\ : LocalMux
    port map (
            O => \N__50152\,
            I => \N__50146\
        );

    \I__11282\ : Odrv4
    port map (
            O => \N__50149\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__11281\ : Odrv4
    port map (
            O => \N__50146\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__11280\ : CascadeMux
    port map (
            O => \N__50141\,
            I => \N__50138\
        );

    \I__11279\ : InMux
    port map (
            O => \N__50138\,
            I => \N__50132\
        );

    \I__11278\ : InMux
    port map (
            O => \N__50137\,
            I => \N__50127\
        );

    \I__11277\ : InMux
    port map (
            O => \N__50136\,
            I => \N__50127\
        );

    \I__11276\ : CascadeMux
    port map (
            O => \N__50135\,
            I => \N__50122\
        );

    \I__11275\ : LocalMux
    port map (
            O => \N__50132\,
            I => \N__50112\
        );

    \I__11274\ : LocalMux
    port map (
            O => \N__50127\,
            I => \N__50112\
        );

    \I__11273\ : CascadeMux
    port map (
            O => \N__50126\,
            I => \N__50108\
        );

    \I__11272\ : InMux
    port map (
            O => \N__50125\,
            I => \N__50092\
        );

    \I__11271\ : InMux
    port map (
            O => \N__50122\,
            I => \N__50068\
        );

    \I__11270\ : InMux
    port map (
            O => \N__50121\,
            I => \N__50068\
        );

    \I__11269\ : InMux
    port map (
            O => \N__50120\,
            I => \N__50068\
        );

    \I__11268\ : InMux
    port map (
            O => \N__50119\,
            I => \N__50068\
        );

    \I__11267\ : InMux
    port map (
            O => \N__50118\,
            I => \N__50068\
        );

    \I__11266\ : InMux
    port map (
            O => \N__50117\,
            I => \N__50068\
        );

    \I__11265\ : Span4Mux_h
    port map (
            O => \N__50112\,
            I => \N__50065\
        );

    \I__11264\ : InMux
    port map (
            O => \N__50111\,
            I => \N__50060\
        );

    \I__11263\ : InMux
    port map (
            O => \N__50108\,
            I => \N__50060\
        );

    \I__11262\ : InMux
    port map (
            O => \N__50107\,
            I => \N__50050\
        );

    \I__11261\ : InMux
    port map (
            O => \N__50106\,
            I => \N__50050\
        );

    \I__11260\ : InMux
    port map (
            O => \N__50105\,
            I => \N__50050\
        );

    \I__11259\ : InMux
    port map (
            O => \N__50104\,
            I => \N__50050\
        );

    \I__11258\ : InMux
    port map (
            O => \N__50103\,
            I => \N__50046\
        );

    \I__11257\ : InMux
    port map (
            O => \N__50102\,
            I => \N__50033\
        );

    \I__11256\ : InMux
    port map (
            O => \N__50101\,
            I => \N__50033\
        );

    \I__11255\ : InMux
    port map (
            O => \N__50100\,
            I => \N__50033\
        );

    \I__11254\ : InMux
    port map (
            O => \N__50099\,
            I => \N__50033\
        );

    \I__11253\ : InMux
    port map (
            O => \N__50098\,
            I => \N__50033\
        );

    \I__11252\ : InMux
    port map (
            O => \N__50097\,
            I => \N__50033\
        );

    \I__11251\ : InMux
    port map (
            O => \N__50096\,
            I => \N__50028\
        );

    \I__11250\ : InMux
    port map (
            O => \N__50095\,
            I => \N__50028\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__50092\,
            I => \N__50025\
        );

    \I__11248\ : InMux
    port map (
            O => \N__50091\,
            I => \N__50022\
        );

    \I__11247\ : InMux
    port map (
            O => \N__50090\,
            I => \N__50004\
        );

    \I__11246\ : InMux
    port map (
            O => \N__50089\,
            I => \N__50004\
        );

    \I__11245\ : InMux
    port map (
            O => \N__50088\,
            I => \N__50004\
        );

    \I__11244\ : InMux
    port map (
            O => \N__50087\,
            I => \N__50004\
        );

    \I__11243\ : InMux
    port map (
            O => \N__50086\,
            I => \N__50004\
        );

    \I__11242\ : InMux
    port map (
            O => \N__50085\,
            I => \N__50004\
        );

    \I__11241\ : InMux
    port map (
            O => \N__50084\,
            I => \N__50004\
        );

    \I__11240\ : InMux
    port map (
            O => \N__50083\,
            I => \N__50004\
        );

    \I__11239\ : InMux
    port map (
            O => \N__50082\,
            I => \N__49999\
        );

    \I__11238\ : InMux
    port map (
            O => \N__50081\,
            I => \N__49999\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__50068\,
            I => \N__49982\
        );

    \I__11236\ : Span4Mux_v
    port map (
            O => \N__50065\,
            I => \N__49973\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__50060\,
            I => \N__49973\
        );

    \I__11234\ : InMux
    port map (
            O => \N__50059\,
            I => \N__49970\
        );

    \I__11233\ : LocalMux
    port map (
            O => \N__50050\,
            I => \N__49967\
        );

    \I__11232\ : InMux
    port map (
            O => \N__50049\,
            I => \N__49964\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__50046\,
            I => \N__49959\
        );

    \I__11230\ : LocalMux
    port map (
            O => \N__50033\,
            I => \N__49959\
        );

    \I__11229\ : LocalMux
    port map (
            O => \N__50028\,
            I => \N__49952\
        );

    \I__11228\ : Span4Mux_h
    port map (
            O => \N__50025\,
            I => \N__49952\
        );

    \I__11227\ : LocalMux
    port map (
            O => \N__50022\,
            I => \N__49952\
        );

    \I__11226\ : CascadeMux
    port map (
            O => \N__50021\,
            I => \N__49937\
        );

    \I__11225\ : LocalMux
    port map (
            O => \N__50004\,
            I => \N__49930\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__49999\,
            I => \N__49930\
        );

    \I__11223\ : InMux
    port map (
            O => \N__49998\,
            I => \N__49923\
        );

    \I__11222\ : InMux
    port map (
            O => \N__49997\,
            I => \N__49923\
        );

    \I__11221\ : InMux
    port map (
            O => \N__49996\,
            I => \N__49923\
        );

    \I__11220\ : InMux
    port map (
            O => \N__49995\,
            I => \N__49912\
        );

    \I__11219\ : InMux
    port map (
            O => \N__49994\,
            I => \N__49912\
        );

    \I__11218\ : InMux
    port map (
            O => \N__49993\,
            I => \N__49912\
        );

    \I__11217\ : InMux
    port map (
            O => \N__49992\,
            I => \N__49912\
        );

    \I__11216\ : InMux
    port map (
            O => \N__49991\,
            I => \N__49912\
        );

    \I__11215\ : InMux
    port map (
            O => \N__49990\,
            I => \N__49899\
        );

    \I__11214\ : InMux
    port map (
            O => \N__49989\,
            I => \N__49899\
        );

    \I__11213\ : InMux
    port map (
            O => \N__49988\,
            I => \N__49899\
        );

    \I__11212\ : InMux
    port map (
            O => \N__49987\,
            I => \N__49899\
        );

    \I__11211\ : InMux
    port map (
            O => \N__49986\,
            I => \N__49899\
        );

    \I__11210\ : InMux
    port map (
            O => \N__49985\,
            I => \N__49899\
        );

    \I__11209\ : Span4Mux_h
    port map (
            O => \N__49982\,
            I => \N__49896\
        );

    \I__11208\ : InMux
    port map (
            O => \N__49981\,
            I => \N__49887\
        );

    \I__11207\ : InMux
    port map (
            O => \N__49980\,
            I => \N__49887\
        );

    \I__11206\ : InMux
    port map (
            O => \N__49979\,
            I => \N__49887\
        );

    \I__11205\ : InMux
    port map (
            O => \N__49978\,
            I => \N__49887\
        );

    \I__11204\ : Span4Mux_h
    port map (
            O => \N__49973\,
            I => \N__49884\
        );

    \I__11203\ : LocalMux
    port map (
            O => \N__49970\,
            I => \N__49881\
        );

    \I__11202\ : Span4Mux_v
    port map (
            O => \N__49967\,
            I => \N__49878\
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__49964\,
            I => \N__49871\
        );

    \I__11200\ : Span4Mux_h
    port map (
            O => \N__49959\,
            I => \N__49871\
        );

    \I__11199\ : Span4Mux_v
    port map (
            O => \N__49952\,
            I => \N__49871\
        );

    \I__11198\ : InMux
    port map (
            O => \N__49951\,
            I => \N__49854\
        );

    \I__11197\ : InMux
    port map (
            O => \N__49950\,
            I => \N__49854\
        );

    \I__11196\ : InMux
    port map (
            O => \N__49949\,
            I => \N__49854\
        );

    \I__11195\ : InMux
    port map (
            O => \N__49948\,
            I => \N__49854\
        );

    \I__11194\ : InMux
    port map (
            O => \N__49947\,
            I => \N__49854\
        );

    \I__11193\ : InMux
    port map (
            O => \N__49946\,
            I => \N__49854\
        );

    \I__11192\ : InMux
    port map (
            O => \N__49945\,
            I => \N__49854\
        );

    \I__11191\ : InMux
    port map (
            O => \N__49944\,
            I => \N__49854\
        );

    \I__11190\ : InMux
    port map (
            O => \N__49943\,
            I => \N__49851\
        );

    \I__11189\ : InMux
    port map (
            O => \N__49942\,
            I => \N__49838\
        );

    \I__11188\ : InMux
    port map (
            O => \N__49941\,
            I => \N__49838\
        );

    \I__11187\ : InMux
    port map (
            O => \N__49940\,
            I => \N__49838\
        );

    \I__11186\ : InMux
    port map (
            O => \N__49937\,
            I => \N__49838\
        );

    \I__11185\ : InMux
    port map (
            O => \N__49936\,
            I => \N__49838\
        );

    \I__11184\ : InMux
    port map (
            O => \N__49935\,
            I => \N__49838\
        );

    \I__11183\ : Span12Mux_h
    port map (
            O => \N__49930\,
            I => \N__49835\
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__49923\,
            I => \N__49824\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__49912\,
            I => \N__49824\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__49899\,
            I => \N__49824\
        );

    \I__11179\ : Sp12to4
    port map (
            O => \N__49896\,
            I => \N__49824\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__49887\,
            I => \N__49824\
        );

    \I__11177\ : Odrv4
    port map (
            O => \N__49884\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11176\ : Odrv4
    port map (
            O => \N__49881\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11175\ : Odrv4
    port map (
            O => \N__49878\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11174\ : Odrv4
    port map (
            O => \N__49871\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11173\ : LocalMux
    port map (
            O => \N__49854\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__49851\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__49838\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11170\ : Odrv12
    port map (
            O => \N__49835\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11169\ : Odrv12
    port map (
            O => \N__49824\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11168\ : CascadeMux
    port map (
            O => \N__49805\,
            I => \N__49801\
        );

    \I__11167\ : InMux
    port map (
            O => \N__49804\,
            I => \N__49796\
        );

    \I__11166\ : InMux
    port map (
            O => \N__49801\,
            I => \N__49796\
        );

    \I__11165\ : LocalMux
    port map (
            O => \N__49796\,
            I => \N__49793\
        );

    \I__11164\ : Span4Mux_v
    port map (
            O => \N__49793\,
            I => \N__49789\
        );

    \I__11163\ : InMux
    port map (
            O => \N__49792\,
            I => \N__49786\
        );

    \I__11162\ : Span4Mux_h
    port map (
            O => \N__49789\,
            I => \N__49782\
        );

    \I__11161\ : LocalMux
    port map (
            O => \N__49786\,
            I => \N__49779\
        );

    \I__11160\ : InMux
    port map (
            O => \N__49785\,
            I => \N__49776\
        );

    \I__11159\ : Odrv4
    port map (
            O => \N__49782\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__11158\ : Odrv12
    port map (
            O => \N__49779\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__49776\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__11156\ : CascadeMux
    port map (
            O => \N__49769\,
            I => \N__49762\
        );

    \I__11155\ : CascadeMux
    port map (
            O => \N__49768\,
            I => \N__49753\
        );

    \I__11154\ : CascadeMux
    port map (
            O => \N__49767\,
            I => \N__49747\
        );

    \I__11153\ : CascadeMux
    port map (
            O => \N__49766\,
            I => \N__49743\
        );

    \I__11152\ : CascadeMux
    port map (
            O => \N__49765\,
            I => \N__49740\
        );

    \I__11151\ : InMux
    port map (
            O => \N__49762\,
            I => \N__49737\
        );

    \I__11150\ : CascadeMux
    port map (
            O => \N__49761\,
            I => \N__49733\
        );

    \I__11149\ : CascadeMux
    port map (
            O => \N__49760\,
            I => \N__49730\
        );

    \I__11148\ : CascadeMux
    port map (
            O => \N__49759\,
            I => \N__49724\
        );

    \I__11147\ : CascadeMux
    port map (
            O => \N__49758\,
            I => \N__49720\
        );

    \I__11146\ : CascadeMux
    port map (
            O => \N__49757\,
            I => \N__49709\
        );

    \I__11145\ : CascadeMux
    port map (
            O => \N__49756\,
            I => \N__49702\
        );

    \I__11144\ : InMux
    port map (
            O => \N__49753\,
            I => \N__49685\
        );

    \I__11143\ : InMux
    port map (
            O => \N__49752\,
            I => \N__49685\
        );

    \I__11142\ : InMux
    port map (
            O => \N__49751\,
            I => \N__49685\
        );

    \I__11141\ : InMux
    port map (
            O => \N__49750\,
            I => \N__49685\
        );

    \I__11140\ : InMux
    port map (
            O => \N__49747\,
            I => \N__49685\
        );

    \I__11139\ : InMux
    port map (
            O => \N__49746\,
            I => \N__49685\
        );

    \I__11138\ : InMux
    port map (
            O => \N__49743\,
            I => \N__49685\
        );

    \I__11137\ : InMux
    port map (
            O => \N__49740\,
            I => \N__49685\
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__49737\,
            I => \N__49682\
        );

    \I__11135\ : InMux
    port map (
            O => \N__49736\,
            I => \N__49667\
        );

    \I__11134\ : InMux
    port map (
            O => \N__49733\,
            I => \N__49667\
        );

    \I__11133\ : InMux
    port map (
            O => \N__49730\,
            I => \N__49667\
        );

    \I__11132\ : InMux
    port map (
            O => \N__49729\,
            I => \N__49667\
        );

    \I__11131\ : InMux
    port map (
            O => \N__49728\,
            I => \N__49667\
        );

    \I__11130\ : InMux
    port map (
            O => \N__49727\,
            I => \N__49667\
        );

    \I__11129\ : InMux
    port map (
            O => \N__49724\,
            I => \N__49667\
        );

    \I__11128\ : InMux
    port map (
            O => \N__49723\,
            I => \N__49662\
        );

    \I__11127\ : InMux
    port map (
            O => \N__49720\,
            I => \N__49662\
        );

    \I__11126\ : InMux
    port map (
            O => \N__49719\,
            I => \N__49651\
        );

    \I__11125\ : InMux
    port map (
            O => \N__49718\,
            I => \N__49651\
        );

    \I__11124\ : InMux
    port map (
            O => \N__49717\,
            I => \N__49651\
        );

    \I__11123\ : InMux
    port map (
            O => \N__49716\,
            I => \N__49651\
        );

    \I__11122\ : InMux
    port map (
            O => \N__49715\,
            I => \N__49651\
        );

    \I__11121\ : InMux
    port map (
            O => \N__49714\,
            I => \N__49640\
        );

    \I__11120\ : InMux
    port map (
            O => \N__49713\,
            I => \N__49640\
        );

    \I__11119\ : InMux
    port map (
            O => \N__49712\,
            I => \N__49640\
        );

    \I__11118\ : InMux
    port map (
            O => \N__49709\,
            I => \N__49640\
        );

    \I__11117\ : CascadeMux
    port map (
            O => \N__49708\,
            I => \N__49636\
        );

    \I__11116\ : CascadeMux
    port map (
            O => \N__49707\,
            I => \N__49631\
        );

    \I__11115\ : CascadeMux
    port map (
            O => \N__49706\,
            I => \N__49628\
        );

    \I__11114\ : CascadeMux
    port map (
            O => \N__49705\,
            I => \N__49625\
        );

    \I__11113\ : InMux
    port map (
            O => \N__49702\,
            I => \N__49609\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__49685\,
            I => \N__49606\
        );

    \I__11111\ : Span4Mux_v
    port map (
            O => \N__49682\,
            I => \N__49597\
        );

    \I__11110\ : LocalMux
    port map (
            O => \N__49667\,
            I => \N__49597\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__49662\,
            I => \N__49597\
        );

    \I__11108\ : LocalMux
    port map (
            O => \N__49651\,
            I => \N__49597\
        );

    \I__11107\ : InMux
    port map (
            O => \N__49650\,
            I => \N__49592\
        );

    \I__11106\ : InMux
    port map (
            O => \N__49649\,
            I => \N__49592\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__49640\,
            I => \N__49589\
        );

    \I__11104\ : InMux
    port map (
            O => \N__49639\,
            I => \N__49586\
        );

    \I__11103\ : InMux
    port map (
            O => \N__49636\,
            I => \N__49583\
        );

    \I__11102\ : InMux
    port map (
            O => \N__49635\,
            I => \N__49572\
        );

    \I__11101\ : InMux
    port map (
            O => \N__49634\,
            I => \N__49572\
        );

    \I__11100\ : InMux
    port map (
            O => \N__49631\,
            I => \N__49572\
        );

    \I__11099\ : InMux
    port map (
            O => \N__49628\,
            I => \N__49572\
        );

    \I__11098\ : InMux
    port map (
            O => \N__49625\,
            I => \N__49572\
        );

    \I__11097\ : InMux
    port map (
            O => \N__49624\,
            I => \N__49569\
        );

    \I__11096\ : InMux
    port map (
            O => \N__49623\,
            I => \N__49564\
        );

    \I__11095\ : InMux
    port map (
            O => \N__49622\,
            I => \N__49564\
        );

    \I__11094\ : CascadeMux
    port map (
            O => \N__49621\,
            I => \N__49535\
        );

    \I__11093\ : CascadeMux
    port map (
            O => \N__49620\,
            I => \N__49531\
        );

    \I__11092\ : CascadeMux
    port map (
            O => \N__49619\,
            I => \N__49527\
        );

    \I__11091\ : CascadeMux
    port map (
            O => \N__49618\,
            I => \N__49523\
        );

    \I__11090\ : CascadeMux
    port map (
            O => \N__49617\,
            I => \N__49519\
        );

    \I__11089\ : CascadeMux
    port map (
            O => \N__49616\,
            I => \N__49515\
        );

    \I__11088\ : CascadeMux
    port map (
            O => \N__49615\,
            I => \N__49511\
        );

    \I__11087\ : CascadeMux
    port map (
            O => \N__49614\,
            I => \N__49496\
        );

    \I__11086\ : CascadeMux
    port map (
            O => \N__49613\,
            I => \N__49492\
        );

    \I__11085\ : CascadeMux
    port map (
            O => \N__49612\,
            I => \N__49488\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__49609\,
            I => \N__49484\
        );

    \I__11083\ : Span4Mux_v
    port map (
            O => \N__49606\,
            I => \N__49477\
        );

    \I__11082\ : Span4Mux_v
    port map (
            O => \N__49597\,
            I => \N__49477\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__49592\,
            I => \N__49477\
        );

    \I__11080\ : Span4Mux_v
    port map (
            O => \N__49589\,
            I => \N__49468\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__49586\,
            I => \N__49468\
        );

    \I__11078\ : LocalMux
    port map (
            O => \N__49583\,
            I => \N__49468\
        );

    \I__11077\ : LocalMux
    port map (
            O => \N__49572\,
            I => \N__49468\
        );

    \I__11076\ : LocalMux
    port map (
            O => \N__49569\,
            I => \N__49463\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__49564\,
            I => \N__49463\
        );

    \I__11074\ : InMux
    port map (
            O => \N__49563\,
            I => \N__49460\
        );

    \I__11073\ : CascadeMux
    port map (
            O => \N__49562\,
            I => \N__49456\
        );

    \I__11072\ : InMux
    port map (
            O => \N__49561\,
            I => \N__49441\
        );

    \I__11071\ : InMux
    port map (
            O => \N__49560\,
            I => \N__49441\
        );

    \I__11070\ : InMux
    port map (
            O => \N__49559\,
            I => \N__49441\
        );

    \I__11069\ : InMux
    port map (
            O => \N__49558\,
            I => \N__49441\
        );

    \I__11068\ : InMux
    port map (
            O => \N__49557\,
            I => \N__49441\
        );

    \I__11067\ : InMux
    port map (
            O => \N__49556\,
            I => \N__49441\
        );

    \I__11066\ : InMux
    port map (
            O => \N__49555\,
            I => \N__49441\
        );

    \I__11065\ : InMux
    port map (
            O => \N__49554\,
            I => \N__49434\
        );

    \I__11064\ : InMux
    port map (
            O => \N__49553\,
            I => \N__49434\
        );

    \I__11063\ : InMux
    port map (
            O => \N__49552\,
            I => \N__49434\
        );

    \I__11062\ : CascadeMux
    port map (
            O => \N__49551\,
            I => \N__49429\
        );

    \I__11061\ : CascadeMux
    port map (
            O => \N__49550\,
            I => \N__49425\
        );

    \I__11060\ : CascadeMux
    port map (
            O => \N__49549\,
            I => \N__49421\
        );

    \I__11059\ : CascadeMux
    port map (
            O => \N__49548\,
            I => \N__49417\
        );

    \I__11058\ : CascadeMux
    port map (
            O => \N__49547\,
            I => \N__49413\
        );

    \I__11057\ : CascadeMux
    port map (
            O => \N__49546\,
            I => \N__49409\
        );

    \I__11056\ : CascadeMux
    port map (
            O => \N__49545\,
            I => \N__49405\
        );

    \I__11055\ : InMux
    port map (
            O => \N__49544\,
            I => \N__49399\
        );

    \I__11054\ : InMux
    port map (
            O => \N__49543\,
            I => \N__49399\
        );

    \I__11053\ : InMux
    port map (
            O => \N__49542\,
            I => \N__49390\
        );

    \I__11052\ : InMux
    port map (
            O => \N__49541\,
            I => \N__49390\
        );

    \I__11051\ : InMux
    port map (
            O => \N__49540\,
            I => \N__49390\
        );

    \I__11050\ : InMux
    port map (
            O => \N__49539\,
            I => \N__49390\
        );

    \I__11049\ : InMux
    port map (
            O => \N__49538\,
            I => \N__49375\
        );

    \I__11048\ : InMux
    port map (
            O => \N__49535\,
            I => \N__49375\
        );

    \I__11047\ : InMux
    port map (
            O => \N__49534\,
            I => \N__49375\
        );

    \I__11046\ : InMux
    port map (
            O => \N__49531\,
            I => \N__49375\
        );

    \I__11045\ : InMux
    port map (
            O => \N__49530\,
            I => \N__49375\
        );

    \I__11044\ : InMux
    port map (
            O => \N__49527\,
            I => \N__49375\
        );

    \I__11043\ : InMux
    port map (
            O => \N__49526\,
            I => \N__49375\
        );

    \I__11042\ : InMux
    port map (
            O => \N__49523\,
            I => \N__49358\
        );

    \I__11041\ : InMux
    port map (
            O => \N__49522\,
            I => \N__49358\
        );

    \I__11040\ : InMux
    port map (
            O => \N__49519\,
            I => \N__49358\
        );

    \I__11039\ : InMux
    port map (
            O => \N__49518\,
            I => \N__49358\
        );

    \I__11038\ : InMux
    port map (
            O => \N__49515\,
            I => \N__49358\
        );

    \I__11037\ : InMux
    port map (
            O => \N__49514\,
            I => \N__49358\
        );

    \I__11036\ : InMux
    port map (
            O => \N__49511\,
            I => \N__49358\
        );

    \I__11035\ : InMux
    port map (
            O => \N__49510\,
            I => \N__49358\
        );

    \I__11034\ : CascadeMux
    port map (
            O => \N__49509\,
            I => \N__49355\
        );

    \I__11033\ : CascadeMux
    port map (
            O => \N__49508\,
            I => \N__49351\
        );

    \I__11032\ : CascadeMux
    port map (
            O => \N__49507\,
            I => \N__49347\
        );

    \I__11031\ : CascadeMux
    port map (
            O => \N__49506\,
            I => \N__49343\
        );

    \I__11030\ : CascadeMux
    port map (
            O => \N__49505\,
            I => \N__49339\
        );

    \I__11029\ : CascadeMux
    port map (
            O => \N__49504\,
            I => \N__49335\
        );

    \I__11028\ : CascadeMux
    port map (
            O => \N__49503\,
            I => \N__49331\
        );

    \I__11027\ : CascadeMux
    port map (
            O => \N__49502\,
            I => \N__49327\
        );

    \I__11026\ : CascadeMux
    port map (
            O => \N__49501\,
            I => \N__49323\
        );

    \I__11025\ : CascadeMux
    port map (
            O => \N__49500\,
            I => \N__49319\
        );

    \I__11024\ : CascadeMux
    port map (
            O => \N__49499\,
            I => \N__49315\
        );

    \I__11023\ : InMux
    port map (
            O => \N__49496\,
            I => \N__49301\
        );

    \I__11022\ : InMux
    port map (
            O => \N__49495\,
            I => \N__49301\
        );

    \I__11021\ : InMux
    port map (
            O => \N__49492\,
            I => \N__49301\
        );

    \I__11020\ : InMux
    port map (
            O => \N__49491\,
            I => \N__49301\
        );

    \I__11019\ : InMux
    port map (
            O => \N__49488\,
            I => \N__49301\
        );

    \I__11018\ : InMux
    port map (
            O => \N__49487\,
            I => \N__49301\
        );

    \I__11017\ : Span12Mux_h
    port map (
            O => \N__49484\,
            I => \N__49298\
        );

    \I__11016\ : Span4Mux_h
    port map (
            O => \N__49477\,
            I => \N__49295\
        );

    \I__11015\ : Span4Mux_h
    port map (
            O => \N__49468\,
            I => \N__49292\
        );

    \I__11014\ : Span4Mux_v
    port map (
            O => \N__49463\,
            I => \N__49287\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__49460\,
            I => \N__49287\
        );

    \I__11012\ : InMux
    port map (
            O => \N__49459\,
            I => \N__49282\
        );

    \I__11011\ : InMux
    port map (
            O => \N__49456\,
            I => \N__49282\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__49441\,
            I => \N__49277\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__49434\,
            I => \N__49277\
        );

    \I__11008\ : InMux
    port map (
            O => \N__49433\,
            I => \N__49260\
        );

    \I__11007\ : InMux
    port map (
            O => \N__49432\,
            I => \N__49260\
        );

    \I__11006\ : InMux
    port map (
            O => \N__49429\,
            I => \N__49260\
        );

    \I__11005\ : InMux
    port map (
            O => \N__49428\,
            I => \N__49260\
        );

    \I__11004\ : InMux
    port map (
            O => \N__49425\,
            I => \N__49260\
        );

    \I__11003\ : InMux
    port map (
            O => \N__49424\,
            I => \N__49260\
        );

    \I__11002\ : InMux
    port map (
            O => \N__49421\,
            I => \N__49260\
        );

    \I__11001\ : InMux
    port map (
            O => \N__49420\,
            I => \N__49260\
        );

    \I__11000\ : InMux
    port map (
            O => \N__49417\,
            I => \N__49243\
        );

    \I__10999\ : InMux
    port map (
            O => \N__49416\,
            I => \N__49243\
        );

    \I__10998\ : InMux
    port map (
            O => \N__49413\,
            I => \N__49243\
        );

    \I__10997\ : InMux
    port map (
            O => \N__49412\,
            I => \N__49243\
        );

    \I__10996\ : InMux
    port map (
            O => \N__49409\,
            I => \N__49243\
        );

    \I__10995\ : InMux
    port map (
            O => \N__49408\,
            I => \N__49243\
        );

    \I__10994\ : InMux
    port map (
            O => \N__49405\,
            I => \N__49243\
        );

    \I__10993\ : InMux
    port map (
            O => \N__49404\,
            I => \N__49243\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__49399\,
            I => \N__49234\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__49390\,
            I => \N__49234\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__49375\,
            I => \N__49234\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__49358\,
            I => \N__49234\
        );

    \I__10988\ : InMux
    port map (
            O => \N__49355\,
            I => \N__49217\
        );

    \I__10987\ : InMux
    port map (
            O => \N__49354\,
            I => \N__49217\
        );

    \I__10986\ : InMux
    port map (
            O => \N__49351\,
            I => \N__49217\
        );

    \I__10985\ : InMux
    port map (
            O => \N__49350\,
            I => \N__49217\
        );

    \I__10984\ : InMux
    port map (
            O => \N__49347\,
            I => \N__49217\
        );

    \I__10983\ : InMux
    port map (
            O => \N__49346\,
            I => \N__49217\
        );

    \I__10982\ : InMux
    port map (
            O => \N__49343\,
            I => \N__49217\
        );

    \I__10981\ : InMux
    port map (
            O => \N__49342\,
            I => \N__49217\
        );

    \I__10980\ : InMux
    port map (
            O => \N__49339\,
            I => \N__49200\
        );

    \I__10979\ : InMux
    port map (
            O => \N__49338\,
            I => \N__49200\
        );

    \I__10978\ : InMux
    port map (
            O => \N__49335\,
            I => \N__49200\
        );

    \I__10977\ : InMux
    port map (
            O => \N__49334\,
            I => \N__49200\
        );

    \I__10976\ : InMux
    port map (
            O => \N__49331\,
            I => \N__49200\
        );

    \I__10975\ : InMux
    port map (
            O => \N__49330\,
            I => \N__49200\
        );

    \I__10974\ : InMux
    port map (
            O => \N__49327\,
            I => \N__49200\
        );

    \I__10973\ : InMux
    port map (
            O => \N__49326\,
            I => \N__49200\
        );

    \I__10972\ : InMux
    port map (
            O => \N__49323\,
            I => \N__49187\
        );

    \I__10971\ : InMux
    port map (
            O => \N__49322\,
            I => \N__49187\
        );

    \I__10970\ : InMux
    port map (
            O => \N__49319\,
            I => \N__49187\
        );

    \I__10969\ : InMux
    port map (
            O => \N__49318\,
            I => \N__49187\
        );

    \I__10968\ : InMux
    port map (
            O => \N__49315\,
            I => \N__49187\
        );

    \I__10967\ : InMux
    port map (
            O => \N__49314\,
            I => \N__49187\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__49301\,
            I => \N__49184\
        );

    \I__10965\ : Odrv12
    port map (
            O => \N__49298\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10964\ : Odrv4
    port map (
            O => \N__49295\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10963\ : Odrv4
    port map (
            O => \N__49292\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10962\ : Odrv4
    port map (
            O => \N__49287\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10961\ : LocalMux
    port map (
            O => \N__49282\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10960\ : Odrv12
    port map (
            O => \N__49277\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__49260\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__49243\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10957\ : Odrv4
    port map (
            O => \N__49234\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10956\ : LocalMux
    port map (
            O => \N__49217\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10955\ : LocalMux
    port map (
            O => \N__49200\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10954\ : LocalMux
    port map (
            O => \N__49187\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10953\ : Odrv4
    port map (
            O => \N__49184\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10952\ : InMux
    port map (
            O => \N__49157\,
            I => \N__49154\
        );

    \I__10951\ : LocalMux
    port map (
            O => \N__49154\,
            I => \N__49151\
        );

    \I__10950\ : Span4Mux_h
    port map (
            O => \N__49151\,
            I => \N__49148\
        );

    \I__10949\ : Odrv4
    port map (
            O => \N__49148\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\
        );

    \I__10948\ : InMux
    port map (
            O => \N__49145\,
            I => \N__49138\
        );

    \I__10947\ : InMux
    port map (
            O => \N__49144\,
            I => \N__49138\
        );

    \I__10946\ : InMux
    port map (
            O => \N__49143\,
            I => \N__49135\
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__49138\,
            I => \N__49130\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__49135\,
            I => \N__49130\
        );

    \I__10943\ : Span4Mux_v
    port map (
            O => \N__49130\,
            I => \N__49125\
        );

    \I__10942\ : CascadeMux
    port map (
            O => \N__49129\,
            I => \N__49122\
        );

    \I__10941\ : CascadeMux
    port map (
            O => \N__49128\,
            I => \N__49119\
        );

    \I__10940\ : Span4Mux_h
    port map (
            O => \N__49125\,
            I => \N__49115\
        );

    \I__10939\ : InMux
    port map (
            O => \N__49122\,
            I => \N__49110\
        );

    \I__10938\ : InMux
    port map (
            O => \N__49119\,
            I => \N__49110\
        );

    \I__10937\ : InMux
    port map (
            O => \N__49118\,
            I => \N__49107\
        );

    \I__10936\ : Span4Mux_h
    port map (
            O => \N__49115\,
            I => \N__49104\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__49110\,
            I => state_3
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__49107\,
            I => state_3
        );

    \I__10933\ : Odrv4
    port map (
            O => \N__49104\,
            I => state_3
        );

    \I__10932\ : IoInMux
    port map (
            O => \N__49097\,
            I => \N__49094\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__49094\,
            I => \N__49091\
        );

    \I__10930\ : Span4Mux_s2_v
    port map (
            O => \N__49091\,
            I => \N__49088\
        );

    \I__10929\ : Span4Mux_v
    port map (
            O => \N__49088\,
            I => \N__49085\
        );

    \I__10928\ : Span4Mux_v
    port map (
            O => \N__49085\,
            I => \N__49080\
        );

    \I__10927\ : InMux
    port map (
            O => \N__49084\,
            I => \N__49075\
        );

    \I__10926\ : InMux
    port map (
            O => \N__49083\,
            I => \N__49075\
        );

    \I__10925\ : Span4Mux_v
    port map (
            O => \N__49080\,
            I => \N__49072\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__49075\,
            I => \N__49069\
        );

    \I__10923\ : Odrv4
    port map (
            O => \N__49072\,
            I => s1_phy_c
        );

    \I__10922\ : Odrv4
    port map (
            O => \N__49069\,
            I => s1_phy_c
        );

    \I__10921\ : InMux
    port map (
            O => \N__49064\,
            I => \N__49058\
        );

    \I__10920\ : InMux
    port map (
            O => \N__49063\,
            I => \N__49055\
        );

    \I__10919\ : InMux
    port map (
            O => \N__49062\,
            I => \N__49052\
        );

    \I__10918\ : InMux
    port map (
            O => \N__49061\,
            I => \N__49049\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__49058\,
            I => \N__49046\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__49055\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__49052\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__10914\ : LocalMux
    port map (
            O => \N__49049\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__10913\ : Odrv4
    port map (
            O => \N__49046\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__10912\ : CascadeMux
    port map (
            O => \N__49037\,
            I => \N__49033\
        );

    \I__10911\ : InMux
    port map (
            O => \N__49036\,
            I => \N__49028\
        );

    \I__10910\ : InMux
    port map (
            O => \N__49033\,
            I => \N__49023\
        );

    \I__10909\ : InMux
    port map (
            O => \N__49032\,
            I => \N__49023\
        );

    \I__10908\ : InMux
    port map (
            O => \N__49031\,
            I => \N__49020\
        );

    \I__10907\ : LocalMux
    port map (
            O => \N__49028\,
            I => \N__49017\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__49023\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__49020\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__10904\ : Odrv4
    port map (
            O => \N__49017\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__10903\ : IoInMux
    port map (
            O => \N__49010\,
            I => \N__49007\
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__49007\,
            I => \N__49004\
        );

    \I__10901\ : Span4Mux_s0_v
    port map (
            O => \N__49004\,
            I => \N__49001\
        );

    \I__10900\ : Span4Mux_h
    port map (
            O => \N__49001\,
            I => \N__48998\
        );

    \I__10899\ : Sp12to4
    port map (
            O => \N__48998\,
            I => \N__48995\
        );

    \I__10898\ : Span12Mux_v
    port map (
            O => \N__48995\,
            I => \N__48992\
        );

    \I__10897\ : Odrv12
    port map (
            O => \N__48992\,
            I => \current_shift_inst.timer_s1.N_163_i\
        );

    \I__10896\ : InMux
    port map (
            O => \N__48989\,
            I => \N__48986\
        );

    \I__10895\ : LocalMux
    port map (
            O => \N__48986\,
            I => \N__48983\
        );

    \I__10894\ : Span4Mux_s2_h
    port map (
            O => \N__48983\,
            I => \N__48979\
        );

    \I__10893\ : InMux
    port map (
            O => \N__48982\,
            I => \N__48976\
        );

    \I__10892\ : Span4Mux_h
    port map (
            O => \N__48979\,
            I => \N__48973\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__48976\,
            I => \N__48968\
        );

    \I__10890\ : Span4Mux_v
    port map (
            O => \N__48973\,
            I => \N__48968\
        );

    \I__10889\ : Odrv4
    port map (
            O => \N__48968\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__10888\ : InMux
    port map (
            O => \N__48965\,
            I => \N__48961\
        );

    \I__10887\ : InMux
    port map (
            O => \N__48964\,
            I => \N__48958\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__48961\,
            I => \N__48955\
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__48958\,
            I => \N__48950\
        );

    \I__10884\ : Span12Mux_s9_v
    port map (
            O => \N__48955\,
            I => \N__48950\
        );

    \I__10883\ : Odrv12
    port map (
            O => \N__48950\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__10882\ : InMux
    port map (
            O => \N__48947\,
            I => \N__48944\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__48944\,
            I => \N__48941\
        );

    \I__10880\ : Span4Mux_s2_h
    port map (
            O => \N__48941\,
            I => \N__48937\
        );

    \I__10879\ : InMux
    port map (
            O => \N__48940\,
            I => \N__48934\
        );

    \I__10878\ : Span4Mux_h
    port map (
            O => \N__48937\,
            I => \N__48931\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__48934\,
            I => \N__48926\
        );

    \I__10876\ : Span4Mux_v
    port map (
            O => \N__48931\,
            I => \N__48926\
        );

    \I__10875\ : Odrv4
    port map (
            O => \N__48926\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__10874\ : InMux
    port map (
            O => \N__48923\,
            I => \N__48920\
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__48920\,
            I => \N__48916\
        );

    \I__10872\ : InMux
    port map (
            O => \N__48919\,
            I => \N__48913\
        );

    \I__10871\ : Span4Mux_v
    port map (
            O => \N__48916\,
            I => \N__48910\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__48913\,
            I => \N__48905\
        );

    \I__10869\ : Span4Mux_h
    port map (
            O => \N__48910\,
            I => \N__48905\
        );

    \I__10868\ : Span4Mux_h
    port map (
            O => \N__48905\,
            I => \N__48902\
        );

    \I__10867\ : Odrv4
    port map (
            O => \N__48902\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__10866\ : CascadeMux
    port map (
            O => \N__48899\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_cascade_\
        );

    \I__10865\ : InMux
    port map (
            O => \N__48896\,
            I => \N__48893\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__48893\,
            I => \N__48890\
        );

    \I__10863\ : Span4Mux_s3_v
    port map (
            O => \N__48890\,
            I => \N__48887\
        );

    \I__10862\ : Odrv4
    port map (
            O => \N__48887\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__10861\ : InMux
    port map (
            O => \N__48884\,
            I => \N__48881\
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__48881\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__10859\ : InMux
    port map (
            O => \N__48878\,
            I => \N__48872\
        );

    \I__10858\ : InMux
    port map (
            O => \N__48877\,
            I => \N__48872\
        );

    \I__10857\ : LocalMux
    port map (
            O => \N__48872\,
            I => \N__48867\
        );

    \I__10856\ : InMux
    port map (
            O => \N__48871\,
            I => \N__48862\
        );

    \I__10855\ : InMux
    port map (
            O => \N__48870\,
            I => \N__48862\
        );

    \I__10854\ : Span4Mux_h
    port map (
            O => \N__48867\,
            I => \N__48859\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__48862\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__10852\ : Odrv4
    port map (
            O => \N__48859\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__10851\ : CascadeMux
    port map (
            O => \N__48854\,
            I => \N__48850\
        );

    \I__10850\ : InMux
    port map (
            O => \N__48853\,
            I => \N__48842\
        );

    \I__10849\ : InMux
    port map (
            O => \N__48850\,
            I => \N__48842\
        );

    \I__10848\ : InMux
    port map (
            O => \N__48849\,
            I => \N__48842\
        );

    \I__10847\ : LocalMux
    port map (
            O => \N__48842\,
            I => \N__48839\
        );

    \I__10846\ : Span4Mux_h
    port map (
            O => \N__48839\,
            I => \N__48836\
        );

    \I__10845\ : Odrv4
    port map (
            O => \N__48836\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__10844\ : ClkMux
    port map (
            O => \N__48833\,
            I => \N__48830\
        );

    \I__10843\ : GlobalMux
    port map (
            O => \N__48830\,
            I => \N__48827\
        );

    \I__10842\ : gio2CtrlBuf
    port map (
            O => \N__48827\,
            I => delay_tr_input_c_g
        );

    \I__10841\ : CEMux
    port map (
            O => \N__48824\,
            I => \N__48821\
        );

    \I__10840\ : LocalMux
    port map (
            O => \N__48821\,
            I => \N__48818\
        );

    \I__10839\ : Span4Mux_v
    port map (
            O => \N__48818\,
            I => \N__48812\
        );

    \I__10838\ : CEMux
    port map (
            O => \N__48817\,
            I => \N__48809\
        );

    \I__10837\ : CEMux
    port map (
            O => \N__48816\,
            I => \N__48806\
        );

    \I__10836\ : CEMux
    port map (
            O => \N__48815\,
            I => \N__48803\
        );

    \I__10835\ : Odrv4
    port map (
            O => \N__48812\,
            I => \current_shift_inst.timer_s1.N_164_i\
        );

    \I__10834\ : LocalMux
    port map (
            O => \N__48809\,
            I => \current_shift_inst.timer_s1.N_164_i\
        );

    \I__10833\ : LocalMux
    port map (
            O => \N__48806\,
            I => \current_shift_inst.timer_s1.N_164_i\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__48803\,
            I => \current_shift_inst.timer_s1.N_164_i\
        );

    \I__10831\ : InMux
    port map (
            O => \N__48794\,
            I => \N__48784\
        );

    \I__10830\ : InMux
    port map (
            O => \N__48793\,
            I => \N__48784\
        );

    \I__10829\ : InMux
    port map (
            O => \N__48792\,
            I => \N__48784\
        );

    \I__10828\ : InMux
    port map (
            O => \N__48791\,
            I => \N__48781\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__48784\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__10826\ : LocalMux
    port map (
            O => \N__48781\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__10825\ : InMux
    port map (
            O => \N__48776\,
            I => \N__48756\
        );

    \I__10824\ : InMux
    port map (
            O => \N__48775\,
            I => \N__48756\
        );

    \I__10823\ : InMux
    port map (
            O => \N__48774\,
            I => \N__48756\
        );

    \I__10822\ : InMux
    port map (
            O => \N__48773\,
            I => \N__48756\
        );

    \I__10821\ : InMux
    port map (
            O => \N__48772\,
            I => \N__48735\
        );

    \I__10820\ : InMux
    port map (
            O => \N__48771\,
            I => \N__48735\
        );

    \I__10819\ : InMux
    port map (
            O => \N__48770\,
            I => \N__48735\
        );

    \I__10818\ : InMux
    port map (
            O => \N__48769\,
            I => \N__48735\
        );

    \I__10817\ : InMux
    port map (
            O => \N__48768\,
            I => \N__48726\
        );

    \I__10816\ : InMux
    port map (
            O => \N__48767\,
            I => \N__48726\
        );

    \I__10815\ : InMux
    port map (
            O => \N__48766\,
            I => \N__48726\
        );

    \I__10814\ : InMux
    port map (
            O => \N__48765\,
            I => \N__48726\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__48756\,
            I => \N__48717\
        );

    \I__10812\ : InMux
    port map (
            O => \N__48755\,
            I => \N__48708\
        );

    \I__10811\ : InMux
    port map (
            O => \N__48754\,
            I => \N__48708\
        );

    \I__10810\ : InMux
    port map (
            O => \N__48753\,
            I => \N__48708\
        );

    \I__10809\ : InMux
    port map (
            O => \N__48752\,
            I => \N__48708\
        );

    \I__10808\ : InMux
    port map (
            O => \N__48751\,
            I => \N__48699\
        );

    \I__10807\ : InMux
    port map (
            O => \N__48750\,
            I => \N__48699\
        );

    \I__10806\ : InMux
    port map (
            O => \N__48749\,
            I => \N__48699\
        );

    \I__10805\ : InMux
    port map (
            O => \N__48748\,
            I => \N__48699\
        );

    \I__10804\ : InMux
    port map (
            O => \N__48747\,
            I => \N__48690\
        );

    \I__10803\ : InMux
    port map (
            O => \N__48746\,
            I => \N__48690\
        );

    \I__10802\ : InMux
    port map (
            O => \N__48745\,
            I => \N__48690\
        );

    \I__10801\ : InMux
    port map (
            O => \N__48744\,
            I => \N__48690\
        );

    \I__10800\ : LocalMux
    port map (
            O => \N__48735\,
            I => \N__48685\
        );

    \I__10799\ : LocalMux
    port map (
            O => \N__48726\,
            I => \N__48685\
        );

    \I__10798\ : InMux
    port map (
            O => \N__48725\,
            I => \N__48680\
        );

    \I__10797\ : InMux
    port map (
            O => \N__48724\,
            I => \N__48680\
        );

    \I__10796\ : InMux
    port map (
            O => \N__48723\,
            I => \N__48671\
        );

    \I__10795\ : InMux
    port map (
            O => \N__48722\,
            I => \N__48671\
        );

    \I__10794\ : InMux
    port map (
            O => \N__48721\,
            I => \N__48671\
        );

    \I__10793\ : InMux
    port map (
            O => \N__48720\,
            I => \N__48671\
        );

    \I__10792\ : Span4Mux_h
    port map (
            O => \N__48717\,
            I => \N__48668\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__48708\,
            I => \N__48659\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__48699\,
            I => \N__48659\
        );

    \I__10789\ : LocalMux
    port map (
            O => \N__48690\,
            I => \N__48659\
        );

    \I__10788\ : Span4Mux_h
    port map (
            O => \N__48685\,
            I => \N__48659\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__48680\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10786\ : LocalMux
    port map (
            O => \N__48671\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10785\ : Odrv4
    port map (
            O => \N__48668\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10784\ : Odrv4
    port map (
            O => \N__48659\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10783\ : InMux
    port map (
            O => \N__48650\,
            I => \N__48647\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__48647\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\
        );

    \I__10781\ : InMux
    port map (
            O => \N__48644\,
            I => \N__48641\
        );

    \I__10780\ : LocalMux
    port map (
            O => \N__48641\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\
        );

    \I__10779\ : CascadeMux
    port map (
            O => \N__48638\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_\
        );

    \I__10778\ : InMux
    port map (
            O => \N__48635\,
            I => \N__48632\
        );

    \I__10777\ : LocalMux
    port map (
            O => \N__48632\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\
        );

    \I__10776\ : InMux
    port map (
            O => \N__48629\,
            I => \N__48626\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__48626\,
            I => \N__48623\
        );

    \I__10774\ : Odrv4
    port map (
            O => \N__48623\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__10773\ : CascadeMux
    port map (
            O => \N__48620\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\
        );

    \I__10772\ : InMux
    port map (
            O => \N__48617\,
            I => \N__48614\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__48614\,
            I => \N__48611\
        );

    \I__10770\ : Odrv12
    port map (
            O => \N__48611\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__10769\ : InMux
    port map (
            O => \N__48608\,
            I => \N__48605\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__48605\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\
        );

    \I__10767\ : InMux
    port map (
            O => \N__48602\,
            I => \N__48599\
        );

    \I__10766\ : LocalMux
    port map (
            O => \N__48599\,
            I => \N__48596\
        );

    \I__10765\ : Odrv4
    port map (
            O => \N__48596\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__10764\ : InMux
    port map (
            O => \N__48593\,
            I => \N__48590\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__48590\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__10762\ : CascadeMux
    port map (
            O => \N__48587\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\
        );

    \I__10761\ : CascadeMux
    port map (
            O => \N__48584\,
            I => \current_shift_inst.PI_CTRL.N_47_cascade_\
        );

    \I__10760\ : InMux
    port map (
            O => \N__48581\,
            I => \N__48578\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__48578\,
            I => \current_shift_inst.PI_CTRL.N_46_21\
        );

    \I__10758\ : CascadeMux
    port map (
            O => \N__48575\,
            I => \N__48572\
        );

    \I__10757\ : InMux
    port map (
            O => \N__48572\,
            I => \N__48569\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__48569\,
            I => \N__48566\
        );

    \I__10755\ : Span4Mux_v
    port map (
            O => \N__48566\,
            I => \N__48563\
        );

    \I__10754\ : Span4Mux_h
    port map (
            O => \N__48563\,
            I => \N__48560\
        );

    \I__10753\ : Odrv4
    port map (
            O => \N__48560\,
            I => \current_shift_inst.PI_CTRL.integrator_1_26\
        );

    \I__10752\ : InMux
    port map (
            O => \N__48557\,
            I => \N__48554\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__48554\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__10750\ : InMux
    port map (
            O => \N__48551\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__10749\ : InMux
    port map (
            O => \N__48548\,
            I => \N__48545\
        );

    \I__10748\ : LocalMux
    port map (
            O => \N__48545\,
            I => \N__48542\
        );

    \I__10747\ : Span12Mux_s6_v
    port map (
            O => \N__48542\,
            I => \N__48539\
        );

    \I__10746\ : Odrv12
    port map (
            O => \N__48539\,
            I => \current_shift_inst.PI_CTRL.integrator_1_27\
        );

    \I__10745\ : InMux
    port map (
            O => \N__48536\,
            I => \N__48533\
        );

    \I__10744\ : LocalMux
    port map (
            O => \N__48533\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__10743\ : InMux
    port map (
            O => \N__48530\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__10742\ : InMux
    port map (
            O => \N__48527\,
            I => \N__48524\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__48524\,
            I => \N__48521\
        );

    \I__10740\ : Span4Mux_h
    port map (
            O => \N__48521\,
            I => \N__48518\
        );

    \I__10739\ : Span4Mux_h
    port map (
            O => \N__48518\,
            I => \N__48515\
        );

    \I__10738\ : Odrv4
    port map (
            O => \N__48515\,
            I => \current_shift_inst.PI_CTRL.integrator_1_28\
        );

    \I__10737\ : InMux
    port map (
            O => \N__48512\,
            I => \N__48509\
        );

    \I__10736\ : LocalMux
    port map (
            O => \N__48509\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__10735\ : InMux
    port map (
            O => \N__48506\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__10734\ : CascadeMux
    port map (
            O => \N__48503\,
            I => \N__48500\
        );

    \I__10733\ : InMux
    port map (
            O => \N__48500\,
            I => \N__48497\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__48497\,
            I => \N__48494\
        );

    \I__10731\ : Span4Mux_h
    port map (
            O => \N__48494\,
            I => \N__48491\
        );

    \I__10730\ : Span4Mux_h
    port map (
            O => \N__48491\,
            I => \N__48488\
        );

    \I__10729\ : Odrv4
    port map (
            O => \N__48488\,
            I => \current_shift_inst.PI_CTRL.integrator_1_29\
        );

    \I__10728\ : InMux
    port map (
            O => \N__48485\,
            I => \N__48482\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__48482\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__10726\ : InMux
    port map (
            O => \N__48479\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__10725\ : InMux
    port map (
            O => \N__48476\,
            I => \N__48473\
        );

    \I__10724\ : LocalMux
    port map (
            O => \N__48473\,
            I => \N__48470\
        );

    \I__10723\ : Span4Mux_h
    port map (
            O => \N__48470\,
            I => \N__48467\
        );

    \I__10722\ : Span4Mux_h
    port map (
            O => \N__48467\,
            I => \N__48464\
        );

    \I__10721\ : Odrv4
    port map (
            O => \N__48464\,
            I => \current_shift_inst.PI_CTRL.integrator_1_30\
        );

    \I__10720\ : InMux
    port map (
            O => \N__48461\,
            I => \N__48458\
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__48458\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__10718\ : InMux
    port map (
            O => \N__48455\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__10717\ : InMux
    port map (
            O => \N__48452\,
            I => \N__48449\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__48449\,
            I => \N__48446\
        );

    \I__10715\ : Span4Mux_v
    port map (
            O => \N__48446\,
            I => \N__48443\
        );

    \I__10714\ : Span4Mux_h
    port map (
            O => \N__48443\,
            I => \N__48440\
        );

    \I__10713\ : Odrv4
    port map (
            O => \N__48440\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30\
        );

    \I__10712\ : CascadeMux
    port map (
            O => \N__48437\,
            I => \N__48434\
        );

    \I__10711\ : InMux
    port map (
            O => \N__48434\,
            I => \N__48431\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__48431\,
            I => \N__48428\
        );

    \I__10709\ : Span4Mux_h
    port map (
            O => \N__48428\,
            I => \N__48425\
        );

    \I__10708\ : Span4Mux_h
    port map (
            O => \N__48425\,
            I => \N__48422\
        );

    \I__10707\ : Odrv4
    port map (
            O => \N__48422\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\
        );

    \I__10706\ : InMux
    port map (
            O => \N__48419\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__10705\ : CascadeMux
    port map (
            O => \N__48416\,
            I => \N__48413\
        );

    \I__10704\ : InMux
    port map (
            O => \N__48413\,
            I => \N__48410\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__48410\,
            I => \N__48407\
        );

    \I__10702\ : Span4Mux_v
    port map (
            O => \N__48407\,
            I => \N__48404\
        );

    \I__10701\ : Span4Mux_h
    port map (
            O => \N__48404\,
            I => \N__48401\
        );

    \I__10700\ : Odrv4
    port map (
            O => \N__48401\,
            I => \current_shift_inst.PI_CTRL.integrator_1_18\
        );

    \I__10699\ : InMux
    port map (
            O => \N__48398\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__10698\ : CascadeMux
    port map (
            O => \N__48395\,
            I => \N__48392\
        );

    \I__10697\ : InMux
    port map (
            O => \N__48392\,
            I => \N__48389\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__48389\,
            I => \N__48386\
        );

    \I__10695\ : Span4Mux_v
    port map (
            O => \N__48386\,
            I => \N__48383\
        );

    \I__10694\ : Span4Mux_h
    port map (
            O => \N__48383\,
            I => \N__48380\
        );

    \I__10693\ : Odrv4
    port map (
            O => \N__48380\,
            I => \current_shift_inst.PI_CTRL.integrator_1_19\
        );

    \I__10692\ : InMux
    port map (
            O => \N__48377\,
            I => \N__48374\
        );

    \I__10691\ : LocalMux
    port map (
            O => \N__48374\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__10690\ : InMux
    port map (
            O => \N__48371\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__10689\ : CascadeMux
    port map (
            O => \N__48368\,
            I => \N__48365\
        );

    \I__10688\ : InMux
    port map (
            O => \N__48365\,
            I => \N__48362\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__48362\,
            I => \N__48359\
        );

    \I__10686\ : Span4Mux_h
    port map (
            O => \N__48359\,
            I => \N__48356\
        );

    \I__10685\ : Span4Mux_h
    port map (
            O => \N__48356\,
            I => \N__48353\
        );

    \I__10684\ : Odrv4
    port map (
            O => \N__48353\,
            I => \current_shift_inst.PI_CTRL.integrator_1_20\
        );

    \I__10683\ : InMux
    port map (
            O => \N__48350\,
            I => \N__48347\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__48347\,
            I => \N__48344\
        );

    \I__10681\ : Span4Mux_h
    port map (
            O => \N__48344\,
            I => \N__48341\
        );

    \I__10680\ : Odrv4
    port map (
            O => \N__48341\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__10679\ : InMux
    port map (
            O => \N__48338\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__10678\ : CascadeMux
    port map (
            O => \N__48335\,
            I => \N__48332\
        );

    \I__10677\ : InMux
    port map (
            O => \N__48332\,
            I => \N__48329\
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__48329\,
            I => \N__48326\
        );

    \I__10675\ : Span4Mux_h
    port map (
            O => \N__48326\,
            I => \N__48323\
        );

    \I__10674\ : Span4Mux_h
    port map (
            O => \N__48323\,
            I => \N__48320\
        );

    \I__10673\ : Odrv4
    port map (
            O => \N__48320\,
            I => \current_shift_inst.PI_CTRL.integrator_1_21\
        );

    \I__10672\ : InMux
    port map (
            O => \N__48317\,
            I => \N__48314\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__48314\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__10670\ : InMux
    port map (
            O => \N__48311\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__10669\ : CascadeMux
    port map (
            O => \N__48308\,
            I => \N__48305\
        );

    \I__10668\ : InMux
    port map (
            O => \N__48305\,
            I => \N__48302\
        );

    \I__10667\ : LocalMux
    port map (
            O => \N__48302\,
            I => \N__48299\
        );

    \I__10666\ : Span4Mux_h
    port map (
            O => \N__48299\,
            I => \N__48296\
        );

    \I__10665\ : Span4Mux_h
    port map (
            O => \N__48296\,
            I => \N__48293\
        );

    \I__10664\ : Odrv4
    port map (
            O => \N__48293\,
            I => \current_shift_inst.PI_CTRL.integrator_1_22\
        );

    \I__10663\ : InMux
    port map (
            O => \N__48290\,
            I => \N__48287\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__48287\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__10661\ : InMux
    port map (
            O => \N__48284\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__10660\ : CascadeMux
    port map (
            O => \N__48281\,
            I => \N__48278\
        );

    \I__10659\ : InMux
    port map (
            O => \N__48278\,
            I => \N__48275\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__48275\,
            I => \N__48272\
        );

    \I__10657\ : Span4Mux_h
    port map (
            O => \N__48272\,
            I => \N__48269\
        );

    \I__10656\ : Span4Mux_h
    port map (
            O => \N__48269\,
            I => \N__48266\
        );

    \I__10655\ : Odrv4
    port map (
            O => \N__48266\,
            I => \current_shift_inst.PI_CTRL.integrator_1_23\
        );

    \I__10654\ : InMux
    port map (
            O => \N__48263\,
            I => \N__48260\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__48260\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__10652\ : InMux
    port map (
            O => \N__48257\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__10651\ : InMux
    port map (
            O => \N__48254\,
            I => \N__48251\
        );

    \I__10650\ : LocalMux
    port map (
            O => \N__48251\,
            I => \N__48248\
        );

    \I__10649\ : Span4Mux_h
    port map (
            O => \N__48248\,
            I => \N__48245\
        );

    \I__10648\ : Span4Mux_h
    port map (
            O => \N__48245\,
            I => \N__48242\
        );

    \I__10647\ : Odrv4
    port map (
            O => \N__48242\,
            I => \current_shift_inst.PI_CTRL.integrator_1_24\
        );

    \I__10646\ : InMux
    port map (
            O => \N__48239\,
            I => \N__48236\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__48236\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__10644\ : InMux
    port map (
            O => \N__48233\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\
        );

    \I__10643\ : InMux
    port map (
            O => \N__48230\,
            I => \N__48227\
        );

    \I__10642\ : LocalMux
    port map (
            O => \N__48227\,
            I => \N__48224\
        );

    \I__10641\ : Span4Mux_h
    port map (
            O => \N__48224\,
            I => \N__48221\
        );

    \I__10640\ : Span4Mux_h
    port map (
            O => \N__48221\,
            I => \N__48218\
        );

    \I__10639\ : Odrv4
    port map (
            O => \N__48218\,
            I => \current_shift_inst.PI_CTRL.integrator_1_25\
        );

    \I__10638\ : InMux
    port map (
            O => \N__48215\,
            I => \N__48212\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__48212\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__10636\ : InMux
    port map (
            O => \N__48209\,
            I => \bfn_17_26_0_\
        );

    \I__10635\ : CascadeMux
    port map (
            O => \N__48206\,
            I => \N__48203\
        );

    \I__10634\ : InMux
    port map (
            O => \N__48203\,
            I => \N__48200\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__48200\,
            I => \N__48197\
        );

    \I__10632\ : Span4Mux_h
    port map (
            O => \N__48197\,
            I => \N__48194\
        );

    \I__10631\ : Span4Mux_h
    port map (
            O => \N__48194\,
            I => \N__48191\
        );

    \I__10630\ : Odrv4
    port map (
            O => \N__48191\,
            I => \current_shift_inst.PI_CTRL.integrator_1_10\
        );

    \I__10629\ : InMux
    port map (
            O => \N__48188\,
            I => \N__48185\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__48185\,
            I => \N__48182\
        );

    \I__10627\ : Span4Mux_v
    port map (
            O => \N__48182\,
            I => \N__48179\
        );

    \I__10626\ : Odrv4
    port map (
            O => \N__48179\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__10625\ : InMux
    port map (
            O => \N__48176\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__10624\ : CascadeMux
    port map (
            O => \N__48173\,
            I => \N__48170\
        );

    \I__10623\ : InMux
    port map (
            O => \N__48170\,
            I => \N__48167\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__48167\,
            I => \N__48164\
        );

    \I__10621\ : Span4Mux_h
    port map (
            O => \N__48164\,
            I => \N__48161\
        );

    \I__10620\ : Span4Mux_h
    port map (
            O => \N__48161\,
            I => \N__48158\
        );

    \I__10619\ : Odrv4
    port map (
            O => \N__48158\,
            I => \current_shift_inst.PI_CTRL.integrator_1_11\
        );

    \I__10618\ : InMux
    port map (
            O => \N__48155\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__10617\ : CascadeMux
    port map (
            O => \N__48152\,
            I => \N__48149\
        );

    \I__10616\ : InMux
    port map (
            O => \N__48149\,
            I => \N__48146\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__48146\,
            I => \N__48143\
        );

    \I__10614\ : Span4Mux_h
    port map (
            O => \N__48143\,
            I => \N__48140\
        );

    \I__10613\ : Span4Mux_h
    port map (
            O => \N__48140\,
            I => \N__48137\
        );

    \I__10612\ : Odrv4
    port map (
            O => \N__48137\,
            I => \current_shift_inst.PI_CTRL.integrator_1_12\
        );

    \I__10611\ : InMux
    port map (
            O => \N__48134\,
            I => \N__48131\
        );

    \I__10610\ : LocalMux
    port map (
            O => \N__48131\,
            I => \N__48128\
        );

    \I__10609\ : Span4Mux_v
    port map (
            O => \N__48128\,
            I => \N__48125\
        );

    \I__10608\ : Odrv4
    port map (
            O => \N__48125\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__10607\ : InMux
    port map (
            O => \N__48122\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__10606\ : CascadeMux
    port map (
            O => \N__48119\,
            I => \N__48116\
        );

    \I__10605\ : InMux
    port map (
            O => \N__48116\,
            I => \N__48113\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__48113\,
            I => \N__48110\
        );

    \I__10603\ : Sp12to4
    port map (
            O => \N__48110\,
            I => \N__48107\
        );

    \I__10602\ : Odrv12
    port map (
            O => \N__48107\,
            I => \current_shift_inst.PI_CTRL.integrator_1_13\
        );

    \I__10601\ : InMux
    port map (
            O => \N__48104\,
            I => \N__48101\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__48101\,
            I => \N__48098\
        );

    \I__10599\ : Span4Mux_s3_v
    port map (
            O => \N__48098\,
            I => \N__48095\
        );

    \I__10598\ : Odrv4
    port map (
            O => \N__48095\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__10597\ : InMux
    port map (
            O => \N__48092\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__10596\ : CascadeMux
    port map (
            O => \N__48089\,
            I => \N__48086\
        );

    \I__10595\ : InMux
    port map (
            O => \N__48086\,
            I => \N__48083\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__48083\,
            I => \N__48080\
        );

    \I__10593\ : Odrv12
    port map (
            O => \N__48080\,
            I => \current_shift_inst.PI_CTRL.integrator_1_14\
        );

    \I__10592\ : InMux
    port map (
            O => \N__48077\,
            I => \N__48074\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__48074\,
            I => \N__48071\
        );

    \I__10590\ : Span4Mux_v
    port map (
            O => \N__48071\,
            I => \N__48068\
        );

    \I__10589\ : Odrv4
    port map (
            O => \N__48068\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__10588\ : InMux
    port map (
            O => \N__48065\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__10587\ : CascadeMux
    port map (
            O => \N__48062\,
            I => \N__48059\
        );

    \I__10586\ : InMux
    port map (
            O => \N__48059\,
            I => \N__48056\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__48056\,
            I => \N__48053\
        );

    \I__10584\ : Sp12to4
    port map (
            O => \N__48053\,
            I => \N__48050\
        );

    \I__10583\ : Odrv12
    port map (
            O => \N__48050\,
            I => \current_shift_inst.PI_CTRL.integrator_1_15\
        );

    \I__10582\ : InMux
    port map (
            O => \N__48047\,
            I => \N__48044\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__48044\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__10580\ : InMux
    port map (
            O => \N__48041\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__10579\ : CascadeMux
    port map (
            O => \N__48038\,
            I => \N__48035\
        );

    \I__10578\ : InMux
    port map (
            O => \N__48035\,
            I => \N__48032\
        );

    \I__10577\ : LocalMux
    port map (
            O => \N__48032\,
            I => \N__48029\
        );

    \I__10576\ : Span4Mux_v
    port map (
            O => \N__48029\,
            I => \N__48026\
        );

    \I__10575\ : Span4Mux_h
    port map (
            O => \N__48026\,
            I => \N__48023\
        );

    \I__10574\ : Odrv4
    port map (
            O => \N__48023\,
            I => \current_shift_inst.PI_CTRL.integrator_1_16\
        );

    \I__10573\ : InMux
    port map (
            O => \N__48020\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\
        );

    \I__10572\ : CascadeMux
    port map (
            O => \N__48017\,
            I => \N__48014\
        );

    \I__10571\ : InMux
    port map (
            O => \N__48014\,
            I => \N__48011\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__48011\,
            I => \N__48008\
        );

    \I__10569\ : Span4Mux_h
    port map (
            O => \N__48008\,
            I => \N__48005\
        );

    \I__10568\ : Span4Mux_h
    port map (
            O => \N__48005\,
            I => \N__48002\
        );

    \I__10567\ : Odrv4
    port map (
            O => \N__48002\,
            I => \current_shift_inst.PI_CTRL.integrator_1_17\
        );

    \I__10566\ : InMux
    port map (
            O => \N__47999\,
            I => \bfn_17_25_0_\
        );

    \I__10565\ : CascadeMux
    port map (
            O => \N__47996\,
            I => \N__47993\
        );

    \I__10564\ : InMux
    port map (
            O => \N__47993\,
            I => \N__47990\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__47990\,
            I => \N__47987\
        );

    \I__10562\ : Span4Mux_h
    port map (
            O => \N__47987\,
            I => \N__47984\
        );

    \I__10561\ : Span4Mux_h
    port map (
            O => \N__47984\,
            I => \N__47981\
        );

    \I__10560\ : Odrv4
    port map (
            O => \N__47981\,
            I => \current_shift_inst.PI_CTRL.integrator_1_2\
        );

    \I__10559\ : InMux
    port map (
            O => \N__47978\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__10558\ : CascadeMux
    port map (
            O => \N__47975\,
            I => \N__47972\
        );

    \I__10557\ : InMux
    port map (
            O => \N__47972\,
            I => \N__47969\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__47969\,
            I => \N__47966\
        );

    \I__10555\ : Span4Mux_h
    port map (
            O => \N__47966\,
            I => \N__47963\
        );

    \I__10554\ : Span4Mux_h
    port map (
            O => \N__47963\,
            I => \N__47960\
        );

    \I__10553\ : Odrv4
    port map (
            O => \N__47960\,
            I => \current_shift_inst.PI_CTRL.integrator_1_3\
        );

    \I__10552\ : InMux
    port map (
            O => \N__47957\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__10551\ : CascadeMux
    port map (
            O => \N__47954\,
            I => \N__47951\
        );

    \I__10550\ : InMux
    port map (
            O => \N__47951\,
            I => \N__47948\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__47948\,
            I => \N__47945\
        );

    \I__10548\ : Span4Mux_h
    port map (
            O => \N__47945\,
            I => \N__47942\
        );

    \I__10547\ : Span4Mux_h
    port map (
            O => \N__47942\,
            I => \N__47939\
        );

    \I__10546\ : Odrv4
    port map (
            O => \N__47939\,
            I => \current_shift_inst.PI_CTRL.integrator_1_4\
        );

    \I__10545\ : InMux
    port map (
            O => \N__47936\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__10544\ : CascadeMux
    port map (
            O => \N__47933\,
            I => \N__47930\
        );

    \I__10543\ : InMux
    port map (
            O => \N__47930\,
            I => \N__47927\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__47927\,
            I => \N__47924\
        );

    \I__10541\ : Span12Mux_v
    port map (
            O => \N__47924\,
            I => \N__47921\
        );

    \I__10540\ : Odrv12
    port map (
            O => \N__47921\,
            I => \current_shift_inst.PI_CTRL.integrator_1_5\
        );

    \I__10539\ : InMux
    port map (
            O => \N__47918\,
            I => \N__47915\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__47915\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__10537\ : InMux
    port map (
            O => \N__47912\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__10536\ : CascadeMux
    port map (
            O => \N__47909\,
            I => \N__47906\
        );

    \I__10535\ : InMux
    port map (
            O => \N__47906\,
            I => \N__47903\
        );

    \I__10534\ : LocalMux
    port map (
            O => \N__47903\,
            I => \N__47900\
        );

    \I__10533\ : Odrv12
    port map (
            O => \N__47900\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__10532\ : InMux
    port map (
            O => \N__47897\,
            I => \N__47894\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__47894\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__10530\ : InMux
    port map (
            O => \N__47891\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__10529\ : CascadeMux
    port map (
            O => \N__47888\,
            I => \N__47885\
        );

    \I__10528\ : InMux
    port map (
            O => \N__47885\,
            I => \N__47882\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__47882\,
            I => \N__47879\
        );

    \I__10526\ : Span12Mux_h
    port map (
            O => \N__47879\,
            I => \N__47876\
        );

    \I__10525\ : Odrv12
    port map (
            O => \N__47876\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__10524\ : InMux
    port map (
            O => \N__47873\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__10523\ : CascadeMux
    port map (
            O => \N__47870\,
            I => \N__47867\
        );

    \I__10522\ : InMux
    port map (
            O => \N__47867\,
            I => \N__47864\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__47864\,
            I => \N__47861\
        );

    \I__10520\ : Odrv12
    port map (
            O => \N__47861\,
            I => \current_shift_inst.PI_CTRL.integrator_1_8\
        );

    \I__10519\ : InMux
    port map (
            O => \N__47858\,
            I => \N__47855\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__47855\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__10517\ : InMux
    port map (
            O => \N__47852\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\
        );

    \I__10516\ : InMux
    port map (
            O => \N__47849\,
            I => \N__47846\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__47846\,
            I => \N__47843\
        );

    \I__10514\ : Span4Mux_h
    port map (
            O => \N__47843\,
            I => \N__47840\
        );

    \I__10513\ : Span4Mux_h
    port map (
            O => \N__47840\,
            I => \N__47837\
        );

    \I__10512\ : Odrv4
    port map (
            O => \N__47837\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__10511\ : InMux
    port map (
            O => \N__47834\,
            I => \bfn_17_24_0_\
        );

    \I__10510\ : InMux
    port map (
            O => \N__47831\,
            I => \N__47828\
        );

    \I__10509\ : LocalMux
    port map (
            O => \N__47828\,
            I => \N__47825\
        );

    \I__10508\ : Span4Mux_h
    port map (
            O => \N__47825\,
            I => \N__47822\
        );

    \I__10507\ : Odrv4
    port map (
            O => \N__47822\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\
        );

    \I__10506\ : InMux
    port map (
            O => \N__47819\,
            I => \bfn_17_22_0_\
        );

    \I__10505\ : InMux
    port map (
            O => \N__47816\,
            I => \N__47813\
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__47813\,
            I => \current_shift_inst.control_input_axb_25\
        );

    \I__10503\ : InMux
    port map (
            O => \N__47810\,
            I => \N__47807\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__47807\,
            I => \N__47804\
        );

    \I__10501\ : Span4Mux_h
    port map (
            O => \N__47804\,
            I => \N__47801\
        );

    \I__10500\ : Odrv4
    port map (
            O => \N__47801\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\
        );

    \I__10499\ : InMux
    port map (
            O => \N__47798\,
            I => \current_shift_inst.control_input_cry_24\
        );

    \I__10498\ : InMux
    port map (
            O => \N__47795\,
            I => \N__47792\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__47792\,
            I => \N__47789\
        );

    \I__10496\ : Span4Mux_v
    port map (
            O => \N__47789\,
            I => \N__47786\
        );

    \I__10495\ : Odrv4
    port map (
            O => \N__47786\,
            I => \current_shift_inst.control_input_axb_26\
        );

    \I__10494\ : InMux
    port map (
            O => \N__47783\,
            I => \N__47780\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__47780\,
            I => \N__47777\
        );

    \I__10492\ : Span4Mux_v
    port map (
            O => \N__47777\,
            I => \N__47774\
        );

    \I__10491\ : Odrv4
    port map (
            O => \N__47774\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\
        );

    \I__10490\ : InMux
    port map (
            O => \N__47771\,
            I => \current_shift_inst.control_input_cry_25\
        );

    \I__10489\ : InMux
    port map (
            O => \N__47768\,
            I => \N__47765\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__47765\,
            I => \current_shift_inst.control_input_axb_27\
        );

    \I__10487\ : InMux
    port map (
            O => \N__47762\,
            I => \N__47759\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__47759\,
            I => \N__47756\
        );

    \I__10485\ : Span4Mux_v
    port map (
            O => \N__47756\,
            I => \N__47753\
        );

    \I__10484\ : Odrv4
    port map (
            O => \N__47753\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\
        );

    \I__10483\ : InMux
    port map (
            O => \N__47750\,
            I => \current_shift_inst.control_input_cry_26\
        );

    \I__10482\ : InMux
    port map (
            O => \N__47747\,
            I => \N__47744\
        );

    \I__10481\ : LocalMux
    port map (
            O => \N__47744\,
            I => \N__47741\
        );

    \I__10480\ : Odrv12
    port map (
            O => \N__47741\,
            I => \current_shift_inst.control_input_axb_28\
        );

    \I__10479\ : InMux
    port map (
            O => \N__47738\,
            I => \N__47735\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__47735\,
            I => \N__47732\
        );

    \I__10477\ : Span4Mux_h
    port map (
            O => \N__47732\,
            I => \N__47729\
        );

    \I__10476\ : Odrv4
    port map (
            O => \N__47729\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\
        );

    \I__10475\ : InMux
    port map (
            O => \N__47726\,
            I => \current_shift_inst.control_input_cry_27\
        );

    \I__10474\ : InMux
    port map (
            O => \N__47723\,
            I => \N__47720\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__47720\,
            I => \N__47717\
        );

    \I__10472\ : Span4Mux_h
    port map (
            O => \N__47717\,
            I => \N__47714\
        );

    \I__10471\ : Odrv4
    port map (
            O => \N__47714\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\
        );

    \I__10470\ : InMux
    port map (
            O => \N__47711\,
            I => \current_shift_inst.control_input_cry_28\
        );

    \I__10469\ : InMux
    port map (
            O => \N__47708\,
            I => \current_shift_inst.control_input_cry_29\
        );

    \I__10468\ : InMux
    port map (
            O => \N__47705\,
            I => \N__47702\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__47702\,
            I => \N__47699\
        );

    \I__10466\ : Span4Mux_h
    port map (
            O => \N__47699\,
            I => \N__47695\
        );

    \I__10465\ : InMux
    port map (
            O => \N__47698\,
            I => \N__47692\
        );

    \I__10464\ : Odrv4
    port map (
            O => \N__47695\,
            I => \current_shift_inst.control_input_31\
        );

    \I__10463\ : LocalMux
    port map (
            O => \N__47692\,
            I => \current_shift_inst.control_input_31\
        );

    \I__10462\ : CascadeMux
    port map (
            O => \N__47687\,
            I => \N__47682\
        );

    \I__10461\ : InMux
    port map (
            O => \N__47686\,
            I => \N__47675\
        );

    \I__10460\ : InMux
    port map (
            O => \N__47685\,
            I => \N__47675\
        );

    \I__10459\ : InMux
    port map (
            O => \N__47682\,
            I => \N__47672\
        );

    \I__10458\ : InMux
    port map (
            O => \N__47681\,
            I => \N__47666\
        );

    \I__10457\ : InMux
    port map (
            O => \N__47680\,
            I => \N__47666\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__47675\,
            I => \N__47656\
        );

    \I__10455\ : LocalMux
    port map (
            O => \N__47672\,
            I => \N__47653\
        );

    \I__10454\ : InMux
    port map (
            O => \N__47671\,
            I => \N__47644\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__47666\,
            I => \N__47641\
        );

    \I__10452\ : InMux
    port map (
            O => \N__47665\,
            I => \N__47636\
        );

    \I__10451\ : InMux
    port map (
            O => \N__47664\,
            I => \N__47636\
        );

    \I__10450\ : InMux
    port map (
            O => \N__47663\,
            I => \N__47625\
        );

    \I__10449\ : InMux
    port map (
            O => \N__47662\,
            I => \N__47625\
        );

    \I__10448\ : InMux
    port map (
            O => \N__47661\,
            I => \N__47625\
        );

    \I__10447\ : InMux
    port map (
            O => \N__47660\,
            I => \N__47625\
        );

    \I__10446\ : InMux
    port map (
            O => \N__47659\,
            I => \N__47625\
        );

    \I__10445\ : Span4Mux_h
    port map (
            O => \N__47656\,
            I => \N__47609\
        );

    \I__10444\ : Span4Mux_h
    port map (
            O => \N__47653\,
            I => \N__47606\
        );

    \I__10443\ : InMux
    port map (
            O => \N__47652\,
            I => \N__47593\
        );

    \I__10442\ : InMux
    port map (
            O => \N__47651\,
            I => \N__47593\
        );

    \I__10441\ : InMux
    port map (
            O => \N__47650\,
            I => \N__47593\
        );

    \I__10440\ : InMux
    port map (
            O => \N__47649\,
            I => \N__47593\
        );

    \I__10439\ : InMux
    port map (
            O => \N__47648\,
            I => \N__47593\
        );

    \I__10438\ : InMux
    port map (
            O => \N__47647\,
            I => \N__47593\
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__47644\,
            I => \N__47584\
        );

    \I__10436\ : Span4Mux_h
    port map (
            O => \N__47641\,
            I => \N__47584\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__47636\,
            I => \N__47584\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__47625\,
            I => \N__47584\
        );

    \I__10433\ : InMux
    port map (
            O => \N__47624\,
            I => \N__47567\
        );

    \I__10432\ : InMux
    port map (
            O => \N__47623\,
            I => \N__47567\
        );

    \I__10431\ : InMux
    port map (
            O => \N__47622\,
            I => \N__47567\
        );

    \I__10430\ : InMux
    port map (
            O => \N__47621\,
            I => \N__47567\
        );

    \I__10429\ : InMux
    port map (
            O => \N__47620\,
            I => \N__47567\
        );

    \I__10428\ : InMux
    port map (
            O => \N__47619\,
            I => \N__47567\
        );

    \I__10427\ : InMux
    port map (
            O => \N__47618\,
            I => \N__47567\
        );

    \I__10426\ : InMux
    port map (
            O => \N__47617\,
            I => \N__47567\
        );

    \I__10425\ : InMux
    port map (
            O => \N__47616\,
            I => \N__47556\
        );

    \I__10424\ : InMux
    port map (
            O => \N__47615\,
            I => \N__47556\
        );

    \I__10423\ : InMux
    port map (
            O => \N__47614\,
            I => \N__47556\
        );

    \I__10422\ : InMux
    port map (
            O => \N__47613\,
            I => \N__47556\
        );

    \I__10421\ : InMux
    port map (
            O => \N__47612\,
            I => \N__47556\
        );

    \I__10420\ : Odrv4
    port map (
            O => \N__47609\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10419\ : Odrv4
    port map (
            O => \N__47606\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__47593\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10417\ : Odrv4
    port map (
            O => \N__47584\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10416\ : LocalMux
    port map (
            O => \N__47567\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__47556\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10414\ : InMux
    port map (
            O => \N__47543\,
            I => \N__47540\
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__47540\,
            I => \current_shift_inst.control_input_axb_29\
        );

    \I__10412\ : CascadeMux
    port map (
            O => \N__47537\,
            I => \N__47534\
        );

    \I__10411\ : InMux
    port map (
            O => \N__47534\,
            I => \N__47531\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__47531\,
            I => \N__47528\
        );

    \I__10409\ : Span4Mux_h
    port map (
            O => \N__47528\,
            I => \N__47525\
        );

    \I__10408\ : Span4Mux_h
    port map (
            O => \N__47525\,
            I => \N__47522\
        );

    \I__10407\ : Odrv4
    port map (
            O => \N__47522\,
            I => \current_shift_inst.PI_CTRL.un1_integrator\
        );

    \I__10406\ : InMux
    port map (
            O => \N__47519\,
            I => \N__47516\
        );

    \I__10405\ : LocalMux
    port map (
            O => \N__47516\,
            I => \current_shift_inst.control_input_axb_17\
        );

    \I__10404\ : InMux
    port map (
            O => \N__47513\,
            I => \N__47510\
        );

    \I__10403\ : LocalMux
    port map (
            O => \N__47510\,
            I => \N__47507\
        );

    \I__10402\ : Span4Mux_h
    port map (
            O => \N__47507\,
            I => \N__47504\
        );

    \I__10401\ : Odrv4
    port map (
            O => \N__47504\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\
        );

    \I__10400\ : InMux
    port map (
            O => \N__47501\,
            I => \current_shift_inst.control_input_cry_16\
        );

    \I__10399\ : InMux
    port map (
            O => \N__47498\,
            I => \N__47495\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__47495\,
            I => \N__47492\
        );

    \I__10397\ : Span4Mux_v
    port map (
            O => \N__47492\,
            I => \N__47489\
        );

    \I__10396\ : Odrv4
    port map (
            O => \N__47489\,
            I => \current_shift_inst.control_input_axb_18\
        );

    \I__10395\ : InMux
    port map (
            O => \N__47486\,
            I => \N__47483\
        );

    \I__10394\ : LocalMux
    port map (
            O => \N__47483\,
            I => \N__47480\
        );

    \I__10393\ : Span4Mux_v
    port map (
            O => \N__47480\,
            I => \N__47477\
        );

    \I__10392\ : Odrv4
    port map (
            O => \N__47477\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\
        );

    \I__10391\ : InMux
    port map (
            O => \N__47474\,
            I => \current_shift_inst.control_input_cry_17\
        );

    \I__10390\ : InMux
    port map (
            O => \N__47471\,
            I => \N__47468\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__47468\,
            I => \N__47465\
        );

    \I__10388\ : Span4Mux_v
    port map (
            O => \N__47465\,
            I => \N__47462\
        );

    \I__10387\ : Odrv4
    port map (
            O => \N__47462\,
            I => \current_shift_inst.control_input_axb_19\
        );

    \I__10386\ : InMux
    port map (
            O => \N__47459\,
            I => \N__47456\
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__47456\,
            I => \N__47453\
        );

    \I__10384\ : Span4Mux_v
    port map (
            O => \N__47453\,
            I => \N__47450\
        );

    \I__10383\ : Odrv4
    port map (
            O => \N__47450\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\
        );

    \I__10382\ : InMux
    port map (
            O => \N__47447\,
            I => \current_shift_inst.control_input_cry_18\
        );

    \I__10381\ : InMux
    port map (
            O => \N__47444\,
            I => \N__47441\
        );

    \I__10380\ : LocalMux
    port map (
            O => \N__47441\,
            I => \current_shift_inst.control_input_axb_20\
        );

    \I__10379\ : InMux
    port map (
            O => \N__47438\,
            I => \N__47435\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__47435\,
            I => \N__47432\
        );

    \I__10377\ : Span4Mux_v
    port map (
            O => \N__47432\,
            I => \N__47429\
        );

    \I__10376\ : Odrv4
    port map (
            O => \N__47429\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\
        );

    \I__10375\ : InMux
    port map (
            O => \N__47426\,
            I => \current_shift_inst.control_input_cry_19\
        );

    \I__10374\ : InMux
    port map (
            O => \N__47423\,
            I => \N__47420\
        );

    \I__10373\ : LocalMux
    port map (
            O => \N__47420\,
            I => \current_shift_inst.control_input_axb_21\
        );

    \I__10372\ : InMux
    port map (
            O => \N__47417\,
            I => \N__47414\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__47414\,
            I => \N__47411\
        );

    \I__10370\ : Span4Mux_h
    port map (
            O => \N__47411\,
            I => \N__47408\
        );

    \I__10369\ : Odrv4
    port map (
            O => \N__47408\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\
        );

    \I__10368\ : InMux
    port map (
            O => \N__47405\,
            I => \current_shift_inst.control_input_cry_20\
        );

    \I__10367\ : InMux
    port map (
            O => \N__47402\,
            I => \N__47399\
        );

    \I__10366\ : LocalMux
    port map (
            O => \N__47399\,
            I => \N__47396\
        );

    \I__10365\ : Odrv4
    port map (
            O => \N__47396\,
            I => \current_shift_inst.control_input_axb_22\
        );

    \I__10364\ : InMux
    port map (
            O => \N__47393\,
            I => \N__47390\
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__47390\,
            I => \N__47387\
        );

    \I__10362\ : Span4Mux_h
    port map (
            O => \N__47387\,
            I => \N__47384\
        );

    \I__10361\ : Odrv4
    port map (
            O => \N__47384\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\
        );

    \I__10360\ : InMux
    port map (
            O => \N__47381\,
            I => \current_shift_inst.control_input_cry_21\
        );

    \I__10359\ : InMux
    port map (
            O => \N__47378\,
            I => \N__47375\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__47375\,
            I => \current_shift_inst.control_input_axb_23\
        );

    \I__10357\ : InMux
    port map (
            O => \N__47372\,
            I => \N__47369\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__47369\,
            I => \N__47366\
        );

    \I__10355\ : Span4Mux_h
    port map (
            O => \N__47366\,
            I => \N__47363\
        );

    \I__10354\ : Odrv4
    port map (
            O => \N__47363\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\
        );

    \I__10353\ : InMux
    port map (
            O => \N__47360\,
            I => \current_shift_inst.control_input_cry_22\
        );

    \I__10352\ : InMux
    port map (
            O => \N__47357\,
            I => \N__47354\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__47354\,
            I => \N__47351\
        );

    \I__10350\ : Span4Mux_v
    port map (
            O => \N__47351\,
            I => \N__47348\
        );

    \I__10349\ : Odrv4
    port map (
            O => \N__47348\,
            I => \current_shift_inst.control_input_axb_24\
        );

    \I__10348\ : InMux
    port map (
            O => \N__47345\,
            I => \N__47342\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__47342\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__10346\ : InMux
    port map (
            O => \N__47339\,
            I => \N__47336\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__47336\,
            I => \N__47333\
        );

    \I__10344\ : Span4Mux_h
    port map (
            O => \N__47333\,
            I => \N__47330\
        );

    \I__10343\ : Odrv4
    port map (
            O => \N__47330\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__10342\ : InMux
    port map (
            O => \N__47327\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__10341\ : InMux
    port map (
            O => \N__47324\,
            I => \N__47321\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__47321\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__10339\ : InMux
    port map (
            O => \N__47318\,
            I => \N__47315\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__47315\,
            I => \N__47312\
        );

    \I__10337\ : Span4Mux_v
    port map (
            O => \N__47312\,
            I => \N__47309\
        );

    \I__10336\ : Odrv4
    port map (
            O => \N__47309\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__10335\ : InMux
    port map (
            O => \N__47306\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__10334\ : InMux
    port map (
            O => \N__47303\,
            I => \N__47300\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__47300\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__10332\ : InMux
    port map (
            O => \N__47297\,
            I => \N__47294\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__47294\,
            I => \N__47291\
        );

    \I__10330\ : Span4Mux_v
    port map (
            O => \N__47291\,
            I => \N__47288\
        );

    \I__10329\ : Odrv4
    port map (
            O => \N__47288\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__10328\ : InMux
    port map (
            O => \N__47285\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__10327\ : InMux
    port map (
            O => \N__47282\,
            I => \N__47279\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__47279\,
            I => \N__47276\
        );

    \I__10325\ : Odrv4
    port map (
            O => \N__47276\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__10324\ : InMux
    port map (
            O => \N__47273\,
            I => \N__47270\
        );

    \I__10323\ : LocalMux
    port map (
            O => \N__47270\,
            I => \N__47267\
        );

    \I__10322\ : Span4Mux_h
    port map (
            O => \N__47267\,
            I => \N__47264\
        );

    \I__10321\ : Odrv4
    port map (
            O => \N__47264\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__10320\ : InMux
    port map (
            O => \N__47261\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__10319\ : InMux
    port map (
            O => \N__47258\,
            I => \N__47255\
        );

    \I__10318\ : LocalMux
    port map (
            O => \N__47255\,
            I => \N__47252\
        );

    \I__10317\ : Odrv4
    port map (
            O => \N__47252\,
            I => \current_shift_inst.control_input_axb_13\
        );

    \I__10316\ : InMux
    port map (
            O => \N__47249\,
            I => \N__47246\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__47246\,
            I => \N__47243\
        );

    \I__10314\ : Span4Mux_h
    port map (
            O => \N__47243\,
            I => \N__47240\
        );

    \I__10313\ : Odrv4
    port map (
            O => \N__47240\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__10312\ : InMux
    port map (
            O => \N__47237\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__10311\ : InMux
    port map (
            O => \N__47234\,
            I => \N__47231\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__47231\,
            I => \N__47228\
        );

    \I__10309\ : Odrv4
    port map (
            O => \N__47228\,
            I => \current_shift_inst.control_input_axb_14\
        );

    \I__10308\ : InMux
    port map (
            O => \N__47225\,
            I => \N__47222\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__47222\,
            I => \N__47219\
        );

    \I__10306\ : Span4Mux_h
    port map (
            O => \N__47219\,
            I => \N__47216\
        );

    \I__10305\ : Odrv4
    port map (
            O => \N__47216\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\
        );

    \I__10304\ : InMux
    port map (
            O => \N__47213\,
            I => \current_shift_inst.control_input_cry_13\
        );

    \I__10303\ : InMux
    port map (
            O => \N__47210\,
            I => \N__47207\
        );

    \I__10302\ : LocalMux
    port map (
            O => \N__47207\,
            I => \current_shift_inst.control_input_axb_15\
        );

    \I__10301\ : InMux
    port map (
            O => \N__47204\,
            I => \N__47201\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__47201\,
            I => \N__47198\
        );

    \I__10299\ : Span4Mux_h
    port map (
            O => \N__47198\,
            I => \N__47195\
        );

    \I__10298\ : Odrv4
    port map (
            O => \N__47195\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\
        );

    \I__10297\ : InMux
    port map (
            O => \N__47192\,
            I => \current_shift_inst.control_input_cry_14\
        );

    \I__10296\ : InMux
    port map (
            O => \N__47189\,
            I => \N__47186\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__47186\,
            I => \N__47183\
        );

    \I__10294\ : Odrv4
    port map (
            O => \N__47183\,
            I => \current_shift_inst.control_input_axb_16\
        );

    \I__10293\ : InMux
    port map (
            O => \N__47180\,
            I => \N__47177\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__47177\,
            I => \N__47174\
        );

    \I__10291\ : Span4Mux_h
    port map (
            O => \N__47174\,
            I => \N__47171\
        );

    \I__10290\ : Odrv4
    port map (
            O => \N__47171\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\
        );

    \I__10289\ : InMux
    port map (
            O => \N__47168\,
            I => \bfn_17_21_0_\
        );

    \I__10288\ : InMux
    port map (
            O => \N__47165\,
            I => \N__47162\
        );

    \I__10287\ : LocalMux
    port map (
            O => \N__47162\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__10286\ : InMux
    port map (
            O => \N__47159\,
            I => \N__47156\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__47156\,
            I => \N__47153\
        );

    \I__10284\ : Span4Mux_h
    port map (
            O => \N__47153\,
            I => \N__47150\
        );

    \I__10283\ : Odrv4
    port map (
            O => \N__47150\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__10282\ : InMux
    port map (
            O => \N__47147\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__10281\ : InMux
    port map (
            O => \N__47144\,
            I => \N__47141\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__47141\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__10279\ : InMux
    port map (
            O => \N__47138\,
            I => \N__47135\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__47135\,
            I => \N__47132\
        );

    \I__10277\ : Span4Mux_v
    port map (
            O => \N__47132\,
            I => \N__47129\
        );

    \I__10276\ : Odrv4
    port map (
            O => \N__47129\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__10275\ : InMux
    port map (
            O => \N__47126\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__10274\ : InMux
    port map (
            O => \N__47123\,
            I => \N__47120\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__47120\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__10272\ : InMux
    port map (
            O => \N__47117\,
            I => \N__47114\
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__47114\,
            I => \N__47111\
        );

    \I__10270\ : Span4Mux_v
    port map (
            O => \N__47111\,
            I => \N__47108\
        );

    \I__10269\ : Odrv4
    port map (
            O => \N__47108\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__10268\ : InMux
    port map (
            O => \N__47105\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__10267\ : InMux
    port map (
            O => \N__47102\,
            I => \N__47099\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__47099\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__10265\ : InMux
    port map (
            O => \N__47096\,
            I => \N__47093\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__47093\,
            I => \N__47090\
        );

    \I__10263\ : Span4Mux_h
    port map (
            O => \N__47090\,
            I => \N__47087\
        );

    \I__10262\ : Odrv4
    port map (
            O => \N__47087\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__10261\ : InMux
    port map (
            O => \N__47084\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__10260\ : InMux
    port map (
            O => \N__47081\,
            I => \N__47078\
        );

    \I__10259\ : LocalMux
    port map (
            O => \N__47078\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__10258\ : InMux
    port map (
            O => \N__47075\,
            I => \N__47072\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__47072\,
            I => \N__47069\
        );

    \I__10256\ : Span4Mux_h
    port map (
            O => \N__47069\,
            I => \N__47066\
        );

    \I__10255\ : Odrv4
    port map (
            O => \N__47066\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__10254\ : InMux
    port map (
            O => \N__47063\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__10253\ : InMux
    port map (
            O => \N__47060\,
            I => \N__47057\
        );

    \I__10252\ : LocalMux
    port map (
            O => \N__47057\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__10251\ : InMux
    port map (
            O => \N__47054\,
            I => \N__47051\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__47051\,
            I => \N__47048\
        );

    \I__10249\ : Span4Mux_h
    port map (
            O => \N__47048\,
            I => \N__47045\
        );

    \I__10248\ : Odrv4
    port map (
            O => \N__47045\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__10247\ : InMux
    port map (
            O => \N__47042\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__10246\ : InMux
    port map (
            O => \N__47039\,
            I => \N__47036\
        );

    \I__10245\ : LocalMux
    port map (
            O => \N__47036\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__10244\ : InMux
    port map (
            O => \N__47033\,
            I => \N__47030\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__47030\,
            I => \N__47027\
        );

    \I__10242\ : Span4Mux_h
    port map (
            O => \N__47027\,
            I => \N__47024\
        );

    \I__10241\ : Odrv4
    port map (
            O => \N__47024\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__10240\ : InMux
    port map (
            O => \N__47021\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__10239\ : InMux
    port map (
            O => \N__47018\,
            I => \N__47015\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__47015\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__10237\ : InMux
    port map (
            O => \N__47012\,
            I => \N__47009\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__47009\,
            I => \N__47006\
        );

    \I__10235\ : Span4Mux_h
    port map (
            O => \N__47006\,
            I => \N__47003\
        );

    \I__10234\ : Odrv4
    port map (
            O => \N__47003\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__10233\ : InMux
    port map (
            O => \N__47000\,
            I => \bfn_17_20_0_\
        );

    \I__10232\ : InMux
    port map (
            O => \N__46997\,
            I => \N__46994\
        );

    \I__10231\ : LocalMux
    port map (
            O => \N__46994\,
            I => \N__46991\
        );

    \I__10230\ : Span12Mux_h
    port map (
            O => \N__46991\,
            I => \N__46988\
        );

    \I__10229\ : Odrv12
    port map (
            O => \N__46988\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__10228\ : InMux
    port map (
            O => \N__46985\,
            I => \N__46982\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__46982\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__10226\ : InMux
    port map (
            O => \N__46979\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__10225\ : CascadeMux
    port map (
            O => \N__46976\,
            I => \N__46973\
        );

    \I__10224\ : InMux
    port map (
            O => \N__46973\,
            I => \N__46970\
        );

    \I__10223\ : LocalMux
    port map (
            O => \N__46970\,
            I => \N__46967\
        );

    \I__10222\ : Odrv12
    port map (
            O => \N__46967\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__10221\ : InMux
    port map (
            O => \N__46964\,
            I => \N__46961\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__46961\,
            I => \N__46958\
        );

    \I__10219\ : Span4Mux_h
    port map (
            O => \N__46958\,
            I => \N__46955\
        );

    \I__10218\ : Odrv4
    port map (
            O => \N__46955\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__10217\ : InMux
    port map (
            O => \N__46952\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__10216\ : InMux
    port map (
            O => \N__46949\,
            I => \N__46946\
        );

    \I__10215\ : LocalMux
    port map (
            O => \N__46946\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__10214\ : InMux
    port map (
            O => \N__46943\,
            I => \N__46940\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__46940\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__10212\ : InMux
    port map (
            O => \N__46937\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__10211\ : CascadeMux
    port map (
            O => \N__46934\,
            I => \N__46931\
        );

    \I__10210\ : InMux
    port map (
            O => \N__46931\,
            I => \N__46928\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__46928\,
            I => \N__46925\
        );

    \I__10208\ : Span4Mux_v
    port map (
            O => \N__46925\,
            I => \N__46922\
        );

    \I__10207\ : Odrv4
    port map (
            O => \N__46922\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__10206\ : InMux
    port map (
            O => \N__46919\,
            I => \N__46916\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__46916\,
            I => \N__46913\
        );

    \I__10204\ : Odrv4
    port map (
            O => \N__46913\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__10203\ : InMux
    port map (
            O => \N__46910\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__10202\ : InMux
    port map (
            O => \N__46907\,
            I => \N__46904\
        );

    \I__10201\ : LocalMux
    port map (
            O => \N__46904\,
            I => \N__46901\
        );

    \I__10200\ : Odrv12
    port map (
            O => \N__46901\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__10199\ : InMux
    port map (
            O => \N__46898\,
            I => \N__46895\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__46895\,
            I => \N__46892\
        );

    \I__10197\ : Sp12to4
    port map (
            O => \N__46892\,
            I => \N__46889\
        );

    \I__10196\ : Odrv12
    port map (
            O => \N__46889\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__10195\ : InMux
    port map (
            O => \N__46886\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__10194\ : CascadeMux
    port map (
            O => \N__46883\,
            I => \N__46880\
        );

    \I__10193\ : InMux
    port map (
            O => \N__46880\,
            I => \N__46877\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__46877\,
            I => \N__46874\
        );

    \I__10191\ : Span4Mux_h
    port map (
            O => \N__46874\,
            I => \N__46871\
        );

    \I__10190\ : Odrv4
    port map (
            O => \N__46871\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__10189\ : InMux
    port map (
            O => \N__46868\,
            I => \N__46865\
        );

    \I__10188\ : LocalMux
    port map (
            O => \N__46865\,
            I => \N__46862\
        );

    \I__10187\ : Odrv4
    port map (
            O => \N__46862\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__10186\ : InMux
    port map (
            O => \N__46859\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__10185\ : InMux
    port map (
            O => \N__46856\,
            I => \N__46853\
        );

    \I__10184\ : LocalMux
    port map (
            O => \N__46853\,
            I => \N__46850\
        );

    \I__10183\ : Span4Mux_h
    port map (
            O => \N__46850\,
            I => \N__46847\
        );

    \I__10182\ : Odrv4
    port map (
            O => \N__46847\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__10181\ : InMux
    port map (
            O => \N__46844\,
            I => \N__46841\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__46841\,
            I => \N__46838\
        );

    \I__10179\ : Odrv4
    port map (
            O => \N__46838\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__10178\ : InMux
    port map (
            O => \N__46835\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__10177\ : InMux
    port map (
            O => \N__46832\,
            I => \N__46829\
        );

    \I__10176\ : LocalMux
    port map (
            O => \N__46829\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__10175\ : CascadeMux
    port map (
            O => \N__46826\,
            I => \N__46821\
        );

    \I__10174\ : InMux
    port map (
            O => \N__46825\,
            I => \N__46818\
        );

    \I__10173\ : InMux
    port map (
            O => \N__46824\,
            I => \N__46815\
        );

    \I__10172\ : InMux
    port map (
            O => \N__46821\,
            I => \N__46812\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__46818\,
            I => \current_shift_inst.N_1619_i\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__46815\,
            I => \current_shift_inst.N_1619_i\
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__46812\,
            I => \current_shift_inst.N_1619_i\
        );

    \I__10168\ : InMux
    port map (
            O => \N__46805\,
            I => \N__46802\
        );

    \I__10167\ : LocalMux
    port map (
            O => \N__46802\,
            I => \N__46799\
        );

    \I__10166\ : Span4Mux_h
    port map (
            O => \N__46799\,
            I => \N__46796\
        );

    \I__10165\ : Odrv4
    port map (
            O => \N__46796\,
            I => \current_shift_inst.control_input_1\
        );

    \I__10164\ : InMux
    port map (
            O => \N__46793\,
            I => \current_shift_inst.un38_control_input_cry_16_s0\
        );

    \I__10163\ : CascadeMux
    port map (
            O => \N__46790\,
            I => \N__46787\
        );

    \I__10162\ : InMux
    port map (
            O => \N__46787\,
            I => \N__46784\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__46784\,
            I => \N__46781\
        );

    \I__10160\ : Span4Mux_h
    port map (
            O => \N__46781\,
            I => \N__46778\
        );

    \I__10159\ : Odrv4
    port map (
            O => \N__46778\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\
        );

    \I__10158\ : InMux
    port map (
            O => \N__46775\,
            I => \N__46772\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__46772\,
            I => \N__46769\
        );

    \I__10156\ : Span4Mux_v
    port map (
            O => \N__46769\,
            I => \N__46766\
        );

    \I__10155\ : Odrv4
    port map (
            O => \N__46766\,
            I => \current_shift_inst.un38_control_input_0_s0_18\
        );

    \I__10154\ : InMux
    port map (
            O => \N__46763\,
            I => \current_shift_inst.un38_control_input_cry_17_s0\
        );

    \I__10153\ : InMux
    port map (
            O => \N__46760\,
            I => \N__46757\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__46757\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\
        );

    \I__10151\ : InMux
    port map (
            O => \N__46754\,
            I => \N__46751\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__46751\,
            I => \current_shift_inst.un38_control_input_0_s0_19\
        );

    \I__10149\ : InMux
    port map (
            O => \N__46748\,
            I => \current_shift_inst.un38_control_input_cry_18_s0\
        );

    \I__10148\ : CascadeMux
    port map (
            O => \N__46745\,
            I => \N__46742\
        );

    \I__10147\ : InMux
    port map (
            O => \N__46742\,
            I => \N__46739\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__46739\,
            I => \N__46736\
        );

    \I__10145\ : Odrv12
    port map (
            O => \N__46736\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__10144\ : InMux
    port map (
            O => \N__46733\,
            I => \N__46730\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__46730\,
            I => \N__46727\
        );

    \I__10142\ : Span4Mux_h
    port map (
            O => \N__46727\,
            I => \N__46724\
        );

    \I__10141\ : Span4Mux_v
    port map (
            O => \N__46724\,
            I => \N__46721\
        );

    \I__10140\ : Odrv4
    port map (
            O => \N__46721\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__10139\ : InMux
    port map (
            O => \N__46718\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__10138\ : InMux
    port map (
            O => \N__46715\,
            I => \N__46712\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__46712\,
            I => \N__46709\
        );

    \I__10136\ : Odrv4
    port map (
            O => \N__46709\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__10135\ : InMux
    port map (
            O => \N__46706\,
            I => \N__46703\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__46703\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__10133\ : InMux
    port map (
            O => \N__46700\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__10132\ : CascadeMux
    port map (
            O => \N__46697\,
            I => \N__46694\
        );

    \I__10131\ : InMux
    port map (
            O => \N__46694\,
            I => \N__46691\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__46691\,
            I => \N__46688\
        );

    \I__10129\ : Span4Mux_h
    port map (
            O => \N__46688\,
            I => \N__46685\
        );

    \I__10128\ : Odrv4
    port map (
            O => \N__46685\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__10127\ : InMux
    port map (
            O => \N__46682\,
            I => \N__46679\
        );

    \I__10126\ : LocalMux
    port map (
            O => \N__46679\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__10125\ : InMux
    port map (
            O => \N__46676\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__10124\ : InMux
    port map (
            O => \N__46673\,
            I => \N__46670\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__46670\,
            I => \N__46667\
        );

    \I__10122\ : Span4Mux_h
    port map (
            O => \N__46667\,
            I => \N__46664\
        );

    \I__10121\ : Odrv4
    port map (
            O => \N__46664\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__10120\ : InMux
    port map (
            O => \N__46661\,
            I => \N__46658\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__46658\,
            I => \N__46655\
        );

    \I__10118\ : Span4Mux_v
    port map (
            O => \N__46655\,
            I => \N__46652\
        );

    \I__10117\ : Odrv4
    port map (
            O => \N__46652\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__10116\ : InMux
    port map (
            O => \N__46649\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__10115\ : CascadeMux
    port map (
            O => \N__46646\,
            I => \N__46643\
        );

    \I__10114\ : InMux
    port map (
            O => \N__46643\,
            I => \N__46640\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__46640\,
            I => \N__46637\
        );

    \I__10112\ : Odrv4
    port map (
            O => \N__46637\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__10111\ : InMux
    port map (
            O => \N__46634\,
            I => \N__46631\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__46631\,
            I => \N__46628\
        );

    \I__10109\ : Span4Mux_v
    port map (
            O => \N__46628\,
            I => \N__46625\
        );

    \I__10108\ : Odrv4
    port map (
            O => \N__46625\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__10107\ : InMux
    port map (
            O => \N__46622\,
            I => \bfn_17_18_0_\
        );

    \I__10106\ : CascadeMux
    port map (
            O => \N__46619\,
            I => \N__46616\
        );

    \I__10105\ : InMux
    port map (
            O => \N__46616\,
            I => \N__46613\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__46613\,
            I => \N__46610\
        );

    \I__10103\ : Span4Mux_h
    port map (
            O => \N__46610\,
            I => \N__46607\
        );

    \I__10102\ : Odrv4
    port map (
            O => \N__46607\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\
        );

    \I__10101\ : InMux
    port map (
            O => \N__46604\,
            I => \N__46601\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__46601\,
            I => \N__46598\
        );

    \I__10099\ : Odrv4
    port map (
            O => \N__46598\,
            I => \current_shift_inst.un38_control_input_0_s0_10\
        );

    \I__10098\ : InMux
    port map (
            O => \N__46595\,
            I => \current_shift_inst.un38_control_input_cry_9_s0\
        );

    \I__10097\ : InMux
    port map (
            O => \N__46592\,
            I => \N__46589\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__46589\,
            I => \N__46586\
        );

    \I__10095\ : Odrv12
    port map (
            O => \N__46586\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\
        );

    \I__10094\ : InMux
    port map (
            O => \N__46583\,
            I => \N__46580\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__46580\,
            I => \N__46577\
        );

    \I__10092\ : Span4Mux_v
    port map (
            O => \N__46577\,
            I => \N__46574\
        );

    \I__10091\ : Odrv4
    port map (
            O => \N__46574\,
            I => \current_shift_inst.un38_control_input_0_s0_11\
        );

    \I__10090\ : InMux
    port map (
            O => \N__46571\,
            I => \current_shift_inst.un38_control_input_cry_10_s0\
        );

    \I__10089\ : CascadeMux
    port map (
            O => \N__46568\,
            I => \N__46565\
        );

    \I__10088\ : InMux
    port map (
            O => \N__46565\,
            I => \N__46562\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__46562\,
            I => \N__46559\
        );

    \I__10086\ : Odrv4
    port map (
            O => \N__46559\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\
        );

    \I__10085\ : InMux
    port map (
            O => \N__46556\,
            I => \N__46553\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__46553\,
            I => \N__46550\
        );

    \I__10083\ : Span4Mux_v
    port map (
            O => \N__46550\,
            I => \N__46547\
        );

    \I__10082\ : Odrv4
    port map (
            O => \N__46547\,
            I => \current_shift_inst.un38_control_input_0_s0_12\
        );

    \I__10081\ : InMux
    port map (
            O => \N__46544\,
            I => \current_shift_inst.un38_control_input_cry_11_s0\
        );

    \I__10080\ : InMux
    port map (
            O => \N__46541\,
            I => \N__46538\
        );

    \I__10079\ : LocalMux
    port map (
            O => \N__46538\,
            I => \N__46535\
        );

    \I__10078\ : Span4Mux_h
    port map (
            O => \N__46535\,
            I => \N__46532\
        );

    \I__10077\ : Odrv4
    port map (
            O => \N__46532\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\
        );

    \I__10076\ : InMux
    port map (
            O => \N__46529\,
            I => \N__46526\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__46526\,
            I => \N__46523\
        );

    \I__10074\ : Span4Mux_v
    port map (
            O => \N__46523\,
            I => \N__46520\
        );

    \I__10073\ : Odrv4
    port map (
            O => \N__46520\,
            I => \current_shift_inst.un38_control_input_0_s0_13\
        );

    \I__10072\ : InMux
    port map (
            O => \N__46517\,
            I => \current_shift_inst.un38_control_input_cry_12_s0\
        );

    \I__10071\ : CascadeMux
    port map (
            O => \N__46514\,
            I => \N__46511\
        );

    \I__10070\ : InMux
    port map (
            O => \N__46511\,
            I => \N__46508\
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__46508\,
            I => \N__46505\
        );

    \I__10068\ : Odrv4
    port map (
            O => \N__46505\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\
        );

    \I__10067\ : InMux
    port map (
            O => \N__46502\,
            I => \N__46499\
        );

    \I__10066\ : LocalMux
    port map (
            O => \N__46499\,
            I => \N__46496\
        );

    \I__10065\ : Span4Mux_v
    port map (
            O => \N__46496\,
            I => \N__46493\
        );

    \I__10064\ : Odrv4
    port map (
            O => \N__46493\,
            I => \current_shift_inst.un38_control_input_0_s0_14\
        );

    \I__10063\ : InMux
    port map (
            O => \N__46490\,
            I => \current_shift_inst.un38_control_input_cry_13_s0\
        );

    \I__10062\ : InMux
    port map (
            O => \N__46487\,
            I => \N__46484\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__46484\,
            I => \N__46481\
        );

    \I__10060\ : Odrv12
    port map (
            O => \N__46481\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\
        );

    \I__10059\ : InMux
    port map (
            O => \N__46478\,
            I => \N__46475\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__46475\,
            I => \N__46472\
        );

    \I__10057\ : Odrv4
    port map (
            O => \N__46472\,
            I => \current_shift_inst.un38_control_input_0_s0_15\
        );

    \I__10056\ : InMux
    port map (
            O => \N__46469\,
            I => \current_shift_inst.un38_control_input_cry_14_s0\
        );

    \I__10055\ : CascadeMux
    port map (
            O => \N__46466\,
            I => \N__46463\
        );

    \I__10054\ : InMux
    port map (
            O => \N__46463\,
            I => \N__46460\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__46460\,
            I => \N__46457\
        );

    \I__10052\ : Span4Mux_h
    port map (
            O => \N__46457\,
            I => \N__46454\
        );

    \I__10051\ : Span4Mux_h
    port map (
            O => \N__46454\,
            I => \N__46451\
        );

    \I__10050\ : Odrv4
    port map (
            O => \N__46451\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\
        );

    \I__10049\ : InMux
    port map (
            O => \N__46448\,
            I => \N__46445\
        );

    \I__10048\ : LocalMux
    port map (
            O => \N__46445\,
            I => \current_shift_inst.un38_control_input_0_s0_16\
        );

    \I__10047\ : InMux
    port map (
            O => \N__46442\,
            I => \bfn_17_17_0_\
        );

    \I__10046\ : InMux
    port map (
            O => \N__46439\,
            I => \N__46436\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__46436\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\
        );

    \I__10044\ : InMux
    port map (
            O => \N__46433\,
            I => \N__46430\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__46430\,
            I => \current_shift_inst.un38_control_input_0_s0_17\
        );

    \I__10042\ : CascadeMux
    port map (
            O => \N__46427\,
            I => \N__46422\
        );

    \I__10041\ : InMux
    port map (
            O => \N__46426\,
            I => \N__46414\
        );

    \I__10040\ : InMux
    port map (
            O => \N__46425\,
            I => \N__46414\
        );

    \I__10039\ : InMux
    port map (
            O => \N__46422\,
            I => \N__46409\
        );

    \I__10038\ : InMux
    port map (
            O => \N__46421\,
            I => \N__46409\
        );

    \I__10037\ : InMux
    port map (
            O => \N__46420\,
            I => \N__46406\
        );

    \I__10036\ : CascadeMux
    port map (
            O => \N__46419\,
            I => \N__46403\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__46414\,
            I => \N__46400\
        );

    \I__10034\ : LocalMux
    port map (
            O => \N__46409\,
            I => \N__46397\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__46406\,
            I => \N__46394\
        );

    \I__10032\ : InMux
    port map (
            O => \N__46403\,
            I => \N__46391\
        );

    \I__10031\ : Span4Mux_h
    port map (
            O => \N__46400\,
            I => \N__46388\
        );

    \I__10030\ : Span4Mux_h
    port map (
            O => \N__46397\,
            I => \N__46381\
        );

    \I__10029\ : Span4Mux_h
    port map (
            O => \N__46394\,
            I => \N__46381\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__46391\,
            I => \N__46381\
        );

    \I__10027\ : Odrv4
    port map (
            O => \N__46388\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__10026\ : Odrv4
    port map (
            O => \N__46381\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__10025\ : CascadeMux
    port map (
            O => \N__46376\,
            I => \N__46373\
        );

    \I__10024\ : InMux
    port map (
            O => \N__46373\,
            I => \N__46370\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__46370\,
            I => \N__46367\
        );

    \I__10022\ : Span4Mux_v
    port map (
            O => \N__46367\,
            I => \N__46364\
        );

    \I__10021\ : Span4Mux_h
    port map (
            O => \N__46364\,
            I => \N__46361\
        );

    \I__10020\ : Odrv4
    port map (
            O => \N__46361\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__10019\ : InMux
    port map (
            O => \N__46358\,
            I => \N__46355\
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__46355\,
            I => \N__46352\
        );

    \I__10017\ : Span4Mux_v
    port map (
            O => \N__46352\,
            I => \N__46349\
        );

    \I__10016\ : Odrv4
    port map (
            O => \N__46349\,
            I => \current_shift_inst.un38_control_input_0_s0_3\
        );

    \I__10015\ : InMux
    port map (
            O => \N__46346\,
            I => \current_shift_inst.un38_control_input_cry_2_s0\
        );

    \I__10014\ : CascadeMux
    port map (
            O => \N__46343\,
            I => \N__46340\
        );

    \I__10013\ : InMux
    port map (
            O => \N__46340\,
            I => \N__46337\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__46337\,
            I => \N__46334\
        );

    \I__10011\ : Span4Mux_h
    port map (
            O => \N__46334\,
            I => \N__46331\
        );

    \I__10010\ : Odrv4
    port map (
            O => \N__46331\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\
        );

    \I__10009\ : InMux
    port map (
            O => \N__46328\,
            I => \N__46325\
        );

    \I__10008\ : LocalMux
    port map (
            O => \N__46325\,
            I => \N__46322\
        );

    \I__10007\ : Span4Mux_v
    port map (
            O => \N__46322\,
            I => \N__46319\
        );

    \I__10006\ : Odrv4
    port map (
            O => \N__46319\,
            I => \current_shift_inst.un38_control_input_0_s0_4\
        );

    \I__10005\ : InMux
    port map (
            O => \N__46316\,
            I => \current_shift_inst.un38_control_input_cry_3_s0\
        );

    \I__10004\ : InMux
    port map (
            O => \N__46313\,
            I => \N__46310\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__46310\,
            I => \N__46307\
        );

    \I__10002\ : Span4Mux_v
    port map (
            O => \N__46307\,
            I => \N__46304\
        );

    \I__10001\ : Odrv4
    port map (
            O => \N__46304\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\
        );

    \I__10000\ : InMux
    port map (
            O => \N__46301\,
            I => \N__46298\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__46298\,
            I => \N__46295\
        );

    \I__9998\ : Sp12to4
    port map (
            O => \N__46295\,
            I => \N__46292\
        );

    \I__9997\ : Odrv12
    port map (
            O => \N__46292\,
            I => \current_shift_inst.un38_control_input_0_s0_5\
        );

    \I__9996\ : InMux
    port map (
            O => \N__46289\,
            I => \current_shift_inst.un38_control_input_cry_4_s0\
        );

    \I__9995\ : CascadeMux
    port map (
            O => \N__46286\,
            I => \N__46283\
        );

    \I__9994\ : InMux
    port map (
            O => \N__46283\,
            I => \N__46280\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__46280\,
            I => \N__46277\
        );

    \I__9992\ : Span4Mux_h
    port map (
            O => \N__46277\,
            I => \N__46274\
        );

    \I__9991\ : Odrv4
    port map (
            O => \N__46274\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\
        );

    \I__9990\ : InMux
    port map (
            O => \N__46271\,
            I => \N__46268\
        );

    \I__9989\ : LocalMux
    port map (
            O => \N__46268\,
            I => \N__46265\
        );

    \I__9988\ : Span4Mux_v
    port map (
            O => \N__46265\,
            I => \N__46262\
        );

    \I__9987\ : Odrv4
    port map (
            O => \N__46262\,
            I => \current_shift_inst.un38_control_input_0_s0_6\
        );

    \I__9986\ : InMux
    port map (
            O => \N__46259\,
            I => \current_shift_inst.un38_control_input_cry_5_s0\
        );

    \I__9985\ : InMux
    port map (
            O => \N__46256\,
            I => \N__46253\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__46253\,
            I => \N__46250\
        );

    \I__9983\ : Span4Mux_v
    port map (
            O => \N__46250\,
            I => \N__46247\
        );

    \I__9982\ : Odrv4
    port map (
            O => \N__46247\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\
        );

    \I__9981\ : InMux
    port map (
            O => \N__46244\,
            I => \N__46241\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__46241\,
            I => \N__46238\
        );

    \I__9979\ : Span4Mux_v
    port map (
            O => \N__46238\,
            I => \N__46235\
        );

    \I__9978\ : Odrv4
    port map (
            O => \N__46235\,
            I => \current_shift_inst.un38_control_input_0_s0_7\
        );

    \I__9977\ : InMux
    port map (
            O => \N__46232\,
            I => \current_shift_inst.un38_control_input_cry_6_s0\
        );

    \I__9976\ : CascadeMux
    port map (
            O => \N__46229\,
            I => \N__46226\
        );

    \I__9975\ : InMux
    port map (
            O => \N__46226\,
            I => \N__46223\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__46223\,
            I => \N__46220\
        );

    \I__9973\ : Span4Mux_h
    port map (
            O => \N__46220\,
            I => \N__46217\
        );

    \I__9972\ : Span4Mux_v
    port map (
            O => \N__46217\,
            I => \N__46214\
        );

    \I__9971\ : Odrv4
    port map (
            O => \N__46214\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\
        );

    \I__9970\ : InMux
    port map (
            O => \N__46211\,
            I => \N__46208\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__46208\,
            I => \N__46205\
        );

    \I__9968\ : Span4Mux_v
    port map (
            O => \N__46205\,
            I => \N__46202\
        );

    \I__9967\ : Odrv4
    port map (
            O => \N__46202\,
            I => \current_shift_inst.un38_control_input_0_s0_8\
        );

    \I__9966\ : InMux
    port map (
            O => \N__46199\,
            I => \bfn_17_16_0_\
        );

    \I__9965\ : InMux
    port map (
            O => \N__46196\,
            I => \N__46193\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__46193\,
            I => \N__46190\
        );

    \I__9963\ : Span4Mux_v
    port map (
            O => \N__46190\,
            I => \N__46187\
        );

    \I__9962\ : Odrv4
    port map (
            O => \N__46187\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\
        );

    \I__9961\ : InMux
    port map (
            O => \N__46184\,
            I => \N__46181\
        );

    \I__9960\ : LocalMux
    port map (
            O => \N__46181\,
            I => \N__46178\
        );

    \I__9959\ : Span4Mux_v
    port map (
            O => \N__46178\,
            I => \N__46175\
        );

    \I__9958\ : Odrv4
    port map (
            O => \N__46175\,
            I => \current_shift_inst.un38_control_input_0_s0_9\
        );

    \I__9957\ : InMux
    port map (
            O => \N__46172\,
            I => \current_shift_inst.un38_control_input_cry_8_s0\
        );

    \I__9956\ : CascadeMux
    port map (
            O => \N__46169\,
            I => \N__46166\
        );

    \I__9955\ : InMux
    port map (
            O => \N__46166\,
            I => \N__46162\
        );

    \I__9954\ : InMux
    port map (
            O => \N__46165\,
            I => \N__46159\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__46162\,
            I => \N__46155\
        );

    \I__9952\ : LocalMux
    port map (
            O => \N__46159\,
            I => \N__46152\
        );

    \I__9951\ : InMux
    port map (
            O => \N__46158\,
            I => \N__46149\
        );

    \I__9950\ : Span4Mux_v
    port map (
            O => \N__46155\,
            I => \N__46146\
        );

    \I__9949\ : Span4Mux_h
    port map (
            O => \N__46152\,
            I => \N__46143\
        );

    \I__9948\ : LocalMux
    port map (
            O => \N__46149\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__9947\ : Odrv4
    port map (
            O => \N__46146\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__9946\ : Odrv4
    port map (
            O => \N__46143\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__9945\ : InMux
    port map (
            O => \N__46136\,
            I => \bfn_17_14_0_\
        );

    \I__9944\ : CascadeMux
    port map (
            O => \N__46133\,
            I => \N__46129\
        );

    \I__9943\ : CascadeMux
    port map (
            O => \N__46132\,
            I => \N__46126\
        );

    \I__9942\ : InMux
    port map (
            O => \N__46129\,
            I => \N__46122\
        );

    \I__9941\ : InMux
    port map (
            O => \N__46126\,
            I => \N__46119\
        );

    \I__9940\ : InMux
    port map (
            O => \N__46125\,
            I => \N__46116\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__46122\,
            I => \N__46113\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__46119\,
            I => \N__46110\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__46116\,
            I => \N__46105\
        );

    \I__9936\ : Span4Mux_v
    port map (
            O => \N__46113\,
            I => \N__46105\
        );

    \I__9935\ : Span4Mux_h
    port map (
            O => \N__46110\,
            I => \N__46102\
        );

    \I__9934\ : Odrv4
    port map (
            O => \N__46105\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__9933\ : Odrv4
    port map (
            O => \N__46102\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__9932\ : InMux
    port map (
            O => \N__46097\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__9931\ : InMux
    port map (
            O => \N__46094\,
            I => \N__46088\
        );

    \I__9930\ : InMux
    port map (
            O => \N__46093\,
            I => \N__46088\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__46088\,
            I => \N__46084\
        );

    \I__9928\ : InMux
    port map (
            O => \N__46087\,
            I => \N__46081\
        );

    \I__9927\ : Span4Mux_h
    port map (
            O => \N__46084\,
            I => \N__46078\
        );

    \I__9926\ : LocalMux
    port map (
            O => \N__46081\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__9925\ : Odrv4
    port map (
            O => \N__46078\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__9924\ : InMux
    port map (
            O => \N__46073\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__9923\ : InMux
    port map (
            O => \N__46070\,
            I => \N__46064\
        );

    \I__9922\ : InMux
    port map (
            O => \N__46069\,
            I => \N__46064\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__46064\,
            I => \N__46060\
        );

    \I__9920\ : InMux
    port map (
            O => \N__46063\,
            I => \N__46057\
        );

    \I__9919\ : Span4Mux_h
    port map (
            O => \N__46060\,
            I => \N__46054\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__46057\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__9917\ : Odrv4
    port map (
            O => \N__46054\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__9916\ : InMux
    port map (
            O => \N__46049\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__9915\ : CascadeMux
    port map (
            O => \N__46046\,
            I => \N__46043\
        );

    \I__9914\ : InMux
    port map (
            O => \N__46043\,
            I => \N__46040\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__46040\,
            I => \N__46037\
        );

    \I__9912\ : Span4Mux_h
    port map (
            O => \N__46037\,
            I => \N__46033\
        );

    \I__9911\ : InMux
    port map (
            O => \N__46036\,
            I => \N__46030\
        );

    \I__9910\ : Span4Mux_h
    port map (
            O => \N__46033\,
            I => \N__46027\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__46030\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__9908\ : Odrv4
    port map (
            O => \N__46027\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__9907\ : InMux
    port map (
            O => \N__46022\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__9906\ : InMux
    port map (
            O => \N__46019\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__9905\ : CascadeMux
    port map (
            O => \N__46016\,
            I => \N__46013\
        );

    \I__9904\ : InMux
    port map (
            O => \N__46013\,
            I => \N__46010\
        );

    \I__9903\ : LocalMux
    port map (
            O => \N__46010\,
            I => \N__46006\
        );

    \I__9902\ : InMux
    port map (
            O => \N__46009\,
            I => \N__46003\
        );

    \I__9901\ : Span4Mux_h
    port map (
            O => \N__46006\,
            I => \N__46000\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__46003\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__9899\ : Odrv4
    port map (
            O => \N__46000\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__9898\ : InMux
    port map (
            O => \N__45995\,
            I => \N__45992\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__45992\,
            I => \N__45989\
        );

    \I__9896\ : Span4Mux_v
    port map (
            O => \N__45989\,
            I => \N__45986\
        );

    \I__9895\ : Odrv4
    port map (
            O => \N__45986\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__9894\ : CascadeMux
    port map (
            O => \N__45983\,
            I => \N__45980\
        );

    \I__9893\ : InMux
    port map (
            O => \N__45980\,
            I => \N__45976\
        );

    \I__9892\ : CascadeMux
    port map (
            O => \N__45979\,
            I => \N__45973\
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__45976\,
            I => \N__45970\
        );

    \I__9890\ : InMux
    port map (
            O => \N__45973\,
            I => \N__45967\
        );

    \I__9889\ : Span4Mux_v
    port map (
            O => \N__45970\,
            I => \N__45962\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__45967\,
            I => \N__45962\
        );

    \I__9887\ : Odrv4
    port map (
            O => \N__45962\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__9886\ : CascadeMux
    port map (
            O => \N__45959\,
            I => \N__45956\
        );

    \I__9885\ : InMux
    port map (
            O => \N__45956\,
            I => \N__45953\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__45953\,
            I => \N__45950\
        );

    \I__9883\ : Span4Mux_h
    port map (
            O => \N__45950\,
            I => \N__45947\
        );

    \I__9882\ : Odrv4
    port map (
            O => \N__45947\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__9881\ : CascadeMux
    port map (
            O => \N__45944\,
            I => \N__45940\
        );

    \I__9880\ : InMux
    port map (
            O => \N__45943\,
            I => \N__45935\
        );

    \I__9879\ : InMux
    port map (
            O => \N__45940\,
            I => \N__45935\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__45935\,
            I => \N__45932\
        );

    \I__9877\ : Span4Mux_v
    port map (
            O => \N__45932\,
            I => \N__45927\
        );

    \I__9876\ : InMux
    port map (
            O => \N__45931\,
            I => \N__45924\
        );

    \I__9875\ : InMux
    port map (
            O => \N__45930\,
            I => \N__45921\
        );

    \I__9874\ : Span4Mux_h
    port map (
            O => \N__45927\,
            I => \N__45916\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__45924\,
            I => \N__45916\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__45921\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__9871\ : Odrv4
    port map (
            O => \N__45916\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__9870\ : InMux
    port map (
            O => \N__45911\,
            I => \N__45905\
        );

    \I__9869\ : InMux
    port map (
            O => \N__45910\,
            I => \N__45905\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__45905\,
            I => \N__45901\
        );

    \I__9867\ : InMux
    port map (
            O => \N__45904\,
            I => \N__45898\
        );

    \I__9866\ : Span4Mux_h
    port map (
            O => \N__45901\,
            I => \N__45895\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__45898\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__9864\ : Odrv4
    port map (
            O => \N__45895\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__9863\ : InMux
    port map (
            O => \N__45890\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__9862\ : CascadeMux
    port map (
            O => \N__45887\,
            I => \N__45884\
        );

    \I__9861\ : InMux
    port map (
            O => \N__45884\,
            I => \N__45879\
        );

    \I__9860\ : InMux
    port map (
            O => \N__45883\,
            I => \N__45876\
        );

    \I__9859\ : InMux
    port map (
            O => \N__45882\,
            I => \N__45873\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__45879\,
            I => \N__45870\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__45876\,
            I => \N__45867\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__45873\,
            I => \N__45862\
        );

    \I__9855\ : Span4Mux_v
    port map (
            O => \N__45870\,
            I => \N__45862\
        );

    \I__9854\ : Span4Mux_h
    port map (
            O => \N__45867\,
            I => \N__45859\
        );

    \I__9853\ : Odrv4
    port map (
            O => \N__45862\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__9852\ : Odrv4
    port map (
            O => \N__45859\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__9851\ : InMux
    port map (
            O => \N__45854\,
            I => \bfn_17_13_0_\
        );

    \I__9850\ : CascadeMux
    port map (
            O => \N__45851\,
            I => \N__45847\
        );

    \I__9849\ : CascadeMux
    port map (
            O => \N__45850\,
            I => \N__45844\
        );

    \I__9848\ : InMux
    port map (
            O => \N__45847\,
            I => \N__45840\
        );

    \I__9847\ : InMux
    port map (
            O => \N__45844\,
            I => \N__45837\
        );

    \I__9846\ : InMux
    port map (
            O => \N__45843\,
            I => \N__45834\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__45840\,
            I => \N__45831\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__45837\,
            I => \N__45828\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__45834\,
            I => \N__45823\
        );

    \I__9842\ : Span4Mux_v
    port map (
            O => \N__45831\,
            I => \N__45823\
        );

    \I__9841\ : Span4Mux_h
    port map (
            O => \N__45828\,
            I => \N__45820\
        );

    \I__9840\ : Odrv4
    port map (
            O => \N__45823\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__9839\ : Odrv4
    port map (
            O => \N__45820\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__9838\ : InMux
    port map (
            O => \N__45815\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__9837\ : CascadeMux
    port map (
            O => \N__45812\,
            I => \N__45809\
        );

    \I__9836\ : InMux
    port map (
            O => \N__45809\,
            I => \N__45805\
        );

    \I__9835\ : InMux
    port map (
            O => \N__45808\,
            I => \N__45802\
        );

    \I__9834\ : LocalMux
    port map (
            O => \N__45805\,
            I => \N__45796\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__45802\,
            I => \N__45796\
        );

    \I__9832\ : InMux
    port map (
            O => \N__45801\,
            I => \N__45793\
        );

    \I__9831\ : Span4Mux_h
    port map (
            O => \N__45796\,
            I => \N__45790\
        );

    \I__9830\ : LocalMux
    port map (
            O => \N__45793\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__9829\ : Odrv4
    port map (
            O => \N__45790\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__9828\ : InMux
    port map (
            O => \N__45785\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__9827\ : InMux
    port map (
            O => \N__45782\,
            I => \N__45776\
        );

    \I__9826\ : InMux
    port map (
            O => \N__45781\,
            I => \N__45776\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__45776\,
            I => \N__45772\
        );

    \I__9824\ : InMux
    port map (
            O => \N__45775\,
            I => \N__45769\
        );

    \I__9823\ : Span4Mux_h
    port map (
            O => \N__45772\,
            I => \N__45766\
        );

    \I__9822\ : LocalMux
    port map (
            O => \N__45769\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__9821\ : Odrv4
    port map (
            O => \N__45766\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__9820\ : InMux
    port map (
            O => \N__45761\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__9819\ : CascadeMux
    port map (
            O => \N__45758\,
            I => \N__45755\
        );

    \I__9818\ : InMux
    port map (
            O => \N__45755\,
            I => \N__45751\
        );

    \I__9817\ : InMux
    port map (
            O => \N__45754\,
            I => \N__45748\
        );

    \I__9816\ : LocalMux
    port map (
            O => \N__45751\,
            I => \N__45742\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__45748\,
            I => \N__45742\
        );

    \I__9814\ : InMux
    port map (
            O => \N__45747\,
            I => \N__45739\
        );

    \I__9813\ : Span4Mux_h
    port map (
            O => \N__45742\,
            I => \N__45736\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__45739\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__9811\ : Odrv4
    port map (
            O => \N__45736\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__9810\ : InMux
    port map (
            O => \N__45731\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__9809\ : CascadeMux
    port map (
            O => \N__45728\,
            I => \N__45724\
        );

    \I__9808\ : CascadeMux
    port map (
            O => \N__45727\,
            I => \N__45721\
        );

    \I__9807\ : InMux
    port map (
            O => \N__45724\,
            I => \N__45716\
        );

    \I__9806\ : InMux
    port map (
            O => \N__45721\,
            I => \N__45716\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__45716\,
            I => \N__45712\
        );

    \I__9804\ : InMux
    port map (
            O => \N__45715\,
            I => \N__45709\
        );

    \I__9803\ : Span4Mux_v
    port map (
            O => \N__45712\,
            I => \N__45706\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__45709\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__9801\ : Odrv4
    port map (
            O => \N__45706\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__9800\ : InMux
    port map (
            O => \N__45701\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__9799\ : CascadeMux
    port map (
            O => \N__45698\,
            I => \N__45695\
        );

    \I__9798\ : InMux
    port map (
            O => \N__45695\,
            I => \N__45691\
        );

    \I__9797\ : InMux
    port map (
            O => \N__45694\,
            I => \N__45688\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__45691\,
            I => \N__45682\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__45688\,
            I => \N__45682\
        );

    \I__9794\ : InMux
    port map (
            O => \N__45687\,
            I => \N__45679\
        );

    \I__9793\ : Span4Mux_v
    port map (
            O => \N__45682\,
            I => \N__45676\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__45679\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__9791\ : Odrv4
    port map (
            O => \N__45676\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__9790\ : InMux
    port map (
            O => \N__45671\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__9789\ : InMux
    port map (
            O => \N__45668\,
            I => \N__45662\
        );

    \I__9788\ : InMux
    port map (
            O => \N__45667\,
            I => \N__45662\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__45662\,
            I => \N__45658\
        );

    \I__9786\ : InMux
    port map (
            O => \N__45661\,
            I => \N__45655\
        );

    \I__9785\ : Span4Mux_h
    port map (
            O => \N__45658\,
            I => \N__45652\
        );

    \I__9784\ : LocalMux
    port map (
            O => \N__45655\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__9783\ : Odrv4
    port map (
            O => \N__45652\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__9782\ : InMux
    port map (
            O => \N__45647\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__9781\ : InMux
    port map (
            O => \N__45644\,
            I => \N__45638\
        );

    \I__9780\ : InMux
    port map (
            O => \N__45643\,
            I => \N__45638\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__45638\,
            I => \N__45634\
        );

    \I__9778\ : InMux
    port map (
            O => \N__45637\,
            I => \N__45631\
        );

    \I__9777\ : Span4Mux_h
    port map (
            O => \N__45634\,
            I => \N__45628\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__45631\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__9775\ : Odrv4
    port map (
            O => \N__45628\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__9774\ : InMux
    port map (
            O => \N__45623\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__9773\ : CascadeMux
    port map (
            O => \N__45620\,
            I => \N__45617\
        );

    \I__9772\ : InMux
    port map (
            O => \N__45617\,
            I => \N__45612\
        );

    \I__9771\ : InMux
    port map (
            O => \N__45616\,
            I => \N__45609\
        );

    \I__9770\ : InMux
    port map (
            O => \N__45615\,
            I => \N__45606\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__45612\,
            I => \N__45603\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__45609\,
            I => \N__45600\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__45606\,
            I => \N__45595\
        );

    \I__9766\ : Span4Mux_v
    port map (
            O => \N__45603\,
            I => \N__45595\
        );

    \I__9765\ : Span4Mux_h
    port map (
            O => \N__45600\,
            I => \N__45592\
        );

    \I__9764\ : Odrv4
    port map (
            O => \N__45595\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__9763\ : Odrv4
    port map (
            O => \N__45592\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__9762\ : InMux
    port map (
            O => \N__45587\,
            I => \bfn_17_12_0_\
        );

    \I__9761\ : CascadeMux
    port map (
            O => \N__45584\,
            I => \N__45580\
        );

    \I__9760\ : CascadeMux
    port map (
            O => \N__45583\,
            I => \N__45577\
        );

    \I__9759\ : InMux
    port map (
            O => \N__45580\,
            I => \N__45574\
        );

    \I__9758\ : InMux
    port map (
            O => \N__45577\,
            I => \N__45571\
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__45574\,
            I => \N__45567\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__45571\,
            I => \N__45564\
        );

    \I__9755\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45561\
        );

    \I__9754\ : Span4Mux_v
    port map (
            O => \N__45567\,
            I => \N__45558\
        );

    \I__9753\ : Span4Mux_h
    port map (
            O => \N__45564\,
            I => \N__45555\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__45561\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__9751\ : Odrv4
    port map (
            O => \N__45558\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__9750\ : Odrv4
    port map (
            O => \N__45555\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__9749\ : InMux
    port map (
            O => \N__45548\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__9748\ : CascadeMux
    port map (
            O => \N__45545\,
            I => \N__45542\
        );

    \I__9747\ : InMux
    port map (
            O => \N__45542\,
            I => \N__45538\
        );

    \I__9746\ : InMux
    port map (
            O => \N__45541\,
            I => \N__45535\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__45538\,
            I => \N__45529\
        );

    \I__9744\ : LocalMux
    port map (
            O => \N__45535\,
            I => \N__45529\
        );

    \I__9743\ : InMux
    port map (
            O => \N__45534\,
            I => \N__45526\
        );

    \I__9742\ : Span4Mux_h
    port map (
            O => \N__45529\,
            I => \N__45523\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__45526\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__9740\ : Odrv4
    port map (
            O => \N__45523\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__9739\ : InMux
    port map (
            O => \N__45518\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__9738\ : InMux
    port map (
            O => \N__45515\,
            I => \N__45509\
        );

    \I__9737\ : InMux
    port map (
            O => \N__45514\,
            I => \N__45509\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__45509\,
            I => \N__45505\
        );

    \I__9735\ : InMux
    port map (
            O => \N__45508\,
            I => \N__45502\
        );

    \I__9734\ : Span4Mux_h
    port map (
            O => \N__45505\,
            I => \N__45499\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__45502\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__9732\ : Odrv4
    port map (
            O => \N__45499\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__9731\ : InMux
    port map (
            O => \N__45494\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__9730\ : InMux
    port map (
            O => \N__45491\,
            I => \N__45485\
        );

    \I__9729\ : InMux
    port map (
            O => \N__45490\,
            I => \N__45485\
        );

    \I__9728\ : LocalMux
    port map (
            O => \N__45485\,
            I => \N__45481\
        );

    \I__9727\ : InMux
    port map (
            O => \N__45484\,
            I => \N__45478\
        );

    \I__9726\ : Span4Mux_h
    port map (
            O => \N__45481\,
            I => \N__45475\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__45478\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__9724\ : Odrv4
    port map (
            O => \N__45475\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__9723\ : InMux
    port map (
            O => \N__45470\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__9722\ : CascadeMux
    port map (
            O => \N__45467\,
            I => \N__45463\
        );

    \I__9721\ : CascadeMux
    port map (
            O => \N__45466\,
            I => \N__45460\
        );

    \I__9720\ : InMux
    port map (
            O => \N__45463\,
            I => \N__45455\
        );

    \I__9719\ : InMux
    port map (
            O => \N__45460\,
            I => \N__45455\
        );

    \I__9718\ : LocalMux
    port map (
            O => \N__45455\,
            I => \N__45451\
        );

    \I__9717\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45448\
        );

    \I__9716\ : Span4Mux_h
    port map (
            O => \N__45451\,
            I => \N__45445\
        );

    \I__9715\ : LocalMux
    port map (
            O => \N__45448\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__9714\ : Odrv4
    port map (
            O => \N__45445\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__9713\ : InMux
    port map (
            O => \N__45440\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__9712\ : CascadeMux
    port map (
            O => \N__45437\,
            I => \N__45433\
        );

    \I__9711\ : CascadeMux
    port map (
            O => \N__45436\,
            I => \N__45430\
        );

    \I__9710\ : InMux
    port map (
            O => \N__45433\,
            I => \N__45425\
        );

    \I__9709\ : InMux
    port map (
            O => \N__45430\,
            I => \N__45425\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__45425\,
            I => \N__45421\
        );

    \I__9707\ : InMux
    port map (
            O => \N__45424\,
            I => \N__45418\
        );

    \I__9706\ : Span4Mux_h
    port map (
            O => \N__45421\,
            I => \N__45415\
        );

    \I__9705\ : LocalMux
    port map (
            O => \N__45418\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__9704\ : Odrv4
    port map (
            O => \N__45415\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__9703\ : InMux
    port map (
            O => \N__45410\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__9702\ : InMux
    port map (
            O => \N__45407\,
            I => \N__45369\
        );

    \I__9701\ : InMux
    port map (
            O => \N__45406\,
            I => \N__45369\
        );

    \I__9700\ : InMux
    port map (
            O => \N__45405\,
            I => \N__45369\
        );

    \I__9699\ : InMux
    port map (
            O => \N__45404\,
            I => \N__45369\
        );

    \I__9698\ : InMux
    port map (
            O => \N__45403\,
            I => \N__45364\
        );

    \I__9697\ : InMux
    port map (
            O => \N__45402\,
            I => \N__45364\
        );

    \I__9696\ : InMux
    port map (
            O => \N__45401\,
            I => \N__45355\
        );

    \I__9695\ : InMux
    port map (
            O => \N__45400\,
            I => \N__45355\
        );

    \I__9694\ : InMux
    port map (
            O => \N__45399\,
            I => \N__45355\
        );

    \I__9693\ : InMux
    port map (
            O => \N__45398\,
            I => \N__45355\
        );

    \I__9692\ : InMux
    port map (
            O => \N__45397\,
            I => \N__45346\
        );

    \I__9691\ : InMux
    port map (
            O => \N__45396\,
            I => \N__45346\
        );

    \I__9690\ : InMux
    port map (
            O => \N__45395\,
            I => \N__45346\
        );

    \I__9689\ : InMux
    port map (
            O => \N__45394\,
            I => \N__45346\
        );

    \I__9688\ : InMux
    port map (
            O => \N__45393\,
            I => \N__45337\
        );

    \I__9687\ : InMux
    port map (
            O => \N__45392\,
            I => \N__45337\
        );

    \I__9686\ : InMux
    port map (
            O => \N__45391\,
            I => \N__45337\
        );

    \I__9685\ : InMux
    port map (
            O => \N__45390\,
            I => \N__45337\
        );

    \I__9684\ : InMux
    port map (
            O => \N__45389\,
            I => \N__45328\
        );

    \I__9683\ : InMux
    port map (
            O => \N__45388\,
            I => \N__45328\
        );

    \I__9682\ : InMux
    port map (
            O => \N__45387\,
            I => \N__45328\
        );

    \I__9681\ : InMux
    port map (
            O => \N__45386\,
            I => \N__45328\
        );

    \I__9680\ : InMux
    port map (
            O => \N__45385\,
            I => \N__45319\
        );

    \I__9679\ : InMux
    port map (
            O => \N__45384\,
            I => \N__45319\
        );

    \I__9678\ : InMux
    port map (
            O => \N__45383\,
            I => \N__45319\
        );

    \I__9677\ : InMux
    port map (
            O => \N__45382\,
            I => \N__45319\
        );

    \I__9676\ : InMux
    port map (
            O => \N__45381\,
            I => \N__45310\
        );

    \I__9675\ : InMux
    port map (
            O => \N__45380\,
            I => \N__45310\
        );

    \I__9674\ : InMux
    port map (
            O => \N__45379\,
            I => \N__45310\
        );

    \I__9673\ : InMux
    port map (
            O => \N__45378\,
            I => \N__45310\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__45369\,
            I => \N__45303\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__45364\,
            I => \N__45303\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__45355\,
            I => \N__45303\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__45346\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__9668\ : LocalMux
    port map (
            O => \N__45337\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__45328\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__45319\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__45310\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__9664\ : Odrv4
    port map (
            O => \N__45303\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__9663\ : InMux
    port map (
            O => \N__45290\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__9662\ : CascadeMux
    port map (
            O => \N__45287\,
            I => \N__45284\
        );

    \I__9661\ : InMux
    port map (
            O => \N__45284\,
            I => \N__45280\
        );

    \I__9660\ : InMux
    port map (
            O => \N__45283\,
            I => \N__45277\
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__45280\,
            I => \N__45274\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__45277\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__9657\ : Odrv12
    port map (
            O => \N__45274\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__9656\ : CEMux
    port map (
            O => \N__45269\,
            I => \N__45264\
        );

    \I__9655\ : CEMux
    port map (
            O => \N__45268\,
            I => \N__45261\
        );

    \I__9654\ : CEMux
    port map (
            O => \N__45267\,
            I => \N__45258\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__45264\,
            I => \N__45255\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__45261\,
            I => \N__45252\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__45258\,
            I => \N__45248\
        );

    \I__9650\ : Span4Mux_v
    port map (
            O => \N__45255\,
            I => \N__45243\
        );

    \I__9649\ : Span4Mux_v
    port map (
            O => \N__45252\,
            I => \N__45243\
        );

    \I__9648\ : CEMux
    port map (
            O => \N__45251\,
            I => \N__45240\
        );

    \I__9647\ : Span4Mux_v
    port map (
            O => \N__45248\,
            I => \N__45233\
        );

    \I__9646\ : Span4Mux_h
    port map (
            O => \N__45243\,
            I => \N__45233\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__45240\,
            I => \N__45233\
        );

    \I__9644\ : Span4Mux_h
    port map (
            O => \N__45233\,
            I => \N__45230\
        );

    \I__9643\ : Odrv4
    port map (
            O => \N__45230\,
            I => \delay_measurement_inst.delay_hc_timer.N_166_i\
        );

    \I__9642\ : InMux
    port map (
            O => \N__45227\,
            I => \N__45224\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__45224\,
            I => \N__45220\
        );

    \I__9640\ : CascadeMux
    port map (
            O => \N__45223\,
            I => \N__45217\
        );

    \I__9639\ : Span4Mux_h
    port map (
            O => \N__45220\,
            I => \N__45213\
        );

    \I__9638\ : InMux
    port map (
            O => \N__45217\,
            I => \N__45210\
        );

    \I__9637\ : InMux
    port map (
            O => \N__45216\,
            I => \N__45207\
        );

    \I__9636\ : Span4Mux_v
    port map (
            O => \N__45213\,
            I => \N__45202\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__45210\,
            I => \N__45202\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__45207\,
            I => \N__45197\
        );

    \I__9633\ : Span4Mux_v
    port map (
            O => \N__45202\,
            I => \N__45197\
        );

    \I__9632\ : Odrv4
    port map (
            O => \N__45197\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__9631\ : InMux
    port map (
            O => \N__45194\,
            I => \bfn_17_11_0_\
        );

    \I__9630\ : InMux
    port map (
            O => \N__45191\,
            I => \N__45187\
        );

    \I__9629\ : CascadeMux
    port map (
            O => \N__45190\,
            I => \N__45184\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__45187\,
            I => \N__45181\
        );

    \I__9627\ : InMux
    port map (
            O => \N__45184\,
            I => \N__45177\
        );

    \I__9626\ : Span4Mux_h
    port map (
            O => \N__45181\,
            I => \N__45174\
        );

    \I__9625\ : InMux
    port map (
            O => \N__45180\,
            I => \N__45171\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__45177\,
            I => \N__45168\
        );

    \I__9623\ : Span4Mux_v
    port map (
            O => \N__45174\,
            I => \N__45165\
        );

    \I__9622\ : LocalMux
    port map (
            O => \N__45171\,
            I => \N__45160\
        );

    \I__9621\ : Span4Mux_v
    port map (
            O => \N__45168\,
            I => \N__45160\
        );

    \I__9620\ : Odrv4
    port map (
            O => \N__45165\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9619\ : Odrv4
    port map (
            O => \N__45160\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9618\ : InMux
    port map (
            O => \N__45155\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__9617\ : InMux
    port map (
            O => \N__45152\,
            I => \N__45146\
        );

    \I__9616\ : InMux
    port map (
            O => \N__45151\,
            I => \N__45146\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__45146\,
            I => \N__45142\
        );

    \I__9614\ : InMux
    port map (
            O => \N__45145\,
            I => \N__45139\
        );

    \I__9613\ : Span4Mux_h
    port map (
            O => \N__45142\,
            I => \N__45136\
        );

    \I__9612\ : LocalMux
    port map (
            O => \N__45139\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__9611\ : Odrv4
    port map (
            O => \N__45136\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__9610\ : InMux
    port map (
            O => \N__45131\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__9609\ : InMux
    port map (
            O => \N__45128\,
            I => \N__45122\
        );

    \I__9608\ : InMux
    port map (
            O => \N__45127\,
            I => \N__45122\
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__45122\,
            I => \N__45118\
        );

    \I__9606\ : InMux
    port map (
            O => \N__45121\,
            I => \N__45115\
        );

    \I__9605\ : Span4Mux_h
    port map (
            O => \N__45118\,
            I => \N__45112\
        );

    \I__9604\ : LocalMux
    port map (
            O => \N__45115\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__9603\ : Odrv4
    port map (
            O => \N__45112\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__9602\ : InMux
    port map (
            O => \N__45107\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__9601\ : CascadeMux
    port map (
            O => \N__45104\,
            I => \N__45100\
        );

    \I__9600\ : CascadeMux
    port map (
            O => \N__45103\,
            I => \N__45097\
        );

    \I__9599\ : InMux
    port map (
            O => \N__45100\,
            I => \N__45092\
        );

    \I__9598\ : InMux
    port map (
            O => \N__45097\,
            I => \N__45092\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__45092\,
            I => \N__45088\
        );

    \I__9596\ : InMux
    port map (
            O => \N__45091\,
            I => \N__45085\
        );

    \I__9595\ : Span4Mux_h
    port map (
            O => \N__45088\,
            I => \N__45082\
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__45085\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__9593\ : Odrv4
    port map (
            O => \N__45082\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__9592\ : InMux
    port map (
            O => \N__45077\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__9591\ : CascadeMux
    port map (
            O => \N__45074\,
            I => \N__45070\
        );

    \I__9590\ : CascadeMux
    port map (
            O => \N__45073\,
            I => \N__45067\
        );

    \I__9589\ : InMux
    port map (
            O => \N__45070\,
            I => \N__45062\
        );

    \I__9588\ : InMux
    port map (
            O => \N__45067\,
            I => \N__45062\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__45062\,
            I => \N__45058\
        );

    \I__9586\ : InMux
    port map (
            O => \N__45061\,
            I => \N__45055\
        );

    \I__9585\ : Span4Mux_h
    port map (
            O => \N__45058\,
            I => \N__45052\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__45055\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__9583\ : Odrv4
    port map (
            O => \N__45052\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__9582\ : InMux
    port map (
            O => \N__45047\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__9581\ : CascadeMux
    port map (
            O => \N__45044\,
            I => \N__45041\
        );

    \I__9580\ : InMux
    port map (
            O => \N__45041\,
            I => \N__45037\
        );

    \I__9579\ : InMux
    port map (
            O => \N__45040\,
            I => \N__45034\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__45037\,
            I => \N__45028\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__45034\,
            I => \N__45028\
        );

    \I__9576\ : InMux
    port map (
            O => \N__45033\,
            I => \N__45025\
        );

    \I__9575\ : Span4Mux_h
    port map (
            O => \N__45028\,
            I => \N__45022\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__45025\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__9573\ : Odrv4
    port map (
            O => \N__45022\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__9572\ : InMux
    port map (
            O => \N__45017\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__9571\ : CascadeMux
    port map (
            O => \N__45014\,
            I => \N__45010\
        );

    \I__9570\ : CascadeMux
    port map (
            O => \N__45013\,
            I => \N__45007\
        );

    \I__9569\ : InMux
    port map (
            O => \N__45010\,
            I => \N__45001\
        );

    \I__9568\ : InMux
    port map (
            O => \N__45007\,
            I => \N__45001\
        );

    \I__9567\ : InMux
    port map (
            O => \N__45006\,
            I => \N__44998\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__45001\,
            I => \N__44995\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__44998\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__9564\ : Odrv12
    port map (
            O => \N__44995\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__9563\ : InMux
    port map (
            O => \N__44990\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__9562\ : CascadeMux
    port map (
            O => \N__44987\,
            I => \N__44983\
        );

    \I__9561\ : CascadeMux
    port map (
            O => \N__44986\,
            I => \N__44980\
        );

    \I__9560\ : InMux
    port map (
            O => \N__44983\,
            I => \N__44974\
        );

    \I__9559\ : InMux
    port map (
            O => \N__44980\,
            I => \N__44974\
        );

    \I__9558\ : InMux
    port map (
            O => \N__44979\,
            I => \N__44971\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__44974\,
            I => \N__44968\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__44971\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__9555\ : Odrv12
    port map (
            O => \N__44968\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__9554\ : InMux
    port map (
            O => \N__44963\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__9553\ : CascadeMux
    port map (
            O => \N__44960\,
            I => \N__44957\
        );

    \I__9552\ : InMux
    port map (
            O => \N__44957\,
            I => \N__44952\
        );

    \I__9551\ : InMux
    port map (
            O => \N__44956\,
            I => \N__44949\
        );

    \I__9550\ : InMux
    port map (
            O => \N__44955\,
            I => \N__44946\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__44952\,
            I => \N__44941\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__44949\,
            I => \N__44941\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__44946\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__9546\ : Odrv12
    port map (
            O => \N__44941\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__9545\ : InMux
    port map (
            O => \N__44936\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__9544\ : CascadeMux
    port map (
            O => \N__44933\,
            I => \N__44930\
        );

    \I__9543\ : InMux
    port map (
            O => \N__44930\,
            I => \N__44925\
        );

    \I__9542\ : InMux
    port map (
            O => \N__44929\,
            I => \N__44922\
        );

    \I__9541\ : InMux
    port map (
            O => \N__44928\,
            I => \N__44919\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__44925\,
            I => \N__44914\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__44922\,
            I => \N__44914\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__44919\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__9537\ : Odrv12
    port map (
            O => \N__44914\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__9536\ : InMux
    port map (
            O => \N__44909\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__9535\ : CascadeMux
    port map (
            O => \N__44906\,
            I => \N__44903\
        );

    \I__9534\ : InMux
    port map (
            O => \N__44903\,
            I => \N__44900\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__44900\,
            I => \N__44895\
        );

    \I__9532\ : InMux
    port map (
            O => \N__44899\,
            I => \N__44892\
        );

    \I__9531\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44889\
        );

    \I__9530\ : Span4Mux_h
    port map (
            O => \N__44895\,
            I => \N__44886\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__44892\,
            I => \N__44883\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__44889\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__9527\ : Odrv4
    port map (
            O => \N__44886\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__9526\ : Odrv12
    port map (
            O => \N__44883\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__9525\ : InMux
    port map (
            O => \N__44876\,
            I => \bfn_17_10_0_\
        );

    \I__9524\ : CascadeMux
    port map (
            O => \N__44873\,
            I => \N__44870\
        );

    \I__9523\ : InMux
    port map (
            O => \N__44870\,
            I => \N__44867\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__44867\,
            I => \N__44862\
        );

    \I__9521\ : InMux
    port map (
            O => \N__44866\,
            I => \N__44859\
        );

    \I__9520\ : InMux
    port map (
            O => \N__44865\,
            I => \N__44856\
        );

    \I__9519\ : Span4Mux_h
    port map (
            O => \N__44862\,
            I => \N__44853\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__44859\,
            I => \N__44850\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__44856\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__9516\ : Odrv4
    port map (
            O => \N__44853\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__9515\ : Odrv12
    port map (
            O => \N__44850\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__9514\ : InMux
    port map (
            O => \N__44843\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__9513\ : InMux
    port map (
            O => \N__44840\,
            I => \N__44833\
        );

    \I__9512\ : InMux
    port map (
            O => \N__44839\,
            I => \N__44833\
        );

    \I__9511\ : InMux
    port map (
            O => \N__44838\,
            I => \N__44830\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__44833\,
            I => \N__44827\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__44830\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__9508\ : Odrv12
    port map (
            O => \N__44827\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__9507\ : InMux
    port map (
            O => \N__44822\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__9506\ : InMux
    port map (
            O => \N__44819\,
            I => \N__44812\
        );

    \I__9505\ : InMux
    port map (
            O => \N__44818\,
            I => \N__44812\
        );

    \I__9504\ : InMux
    port map (
            O => \N__44817\,
            I => \N__44809\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__44812\,
            I => \N__44806\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__44809\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__9501\ : Odrv12
    port map (
            O => \N__44806\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__9500\ : InMux
    port map (
            O => \N__44801\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__9499\ : CascadeMux
    port map (
            O => \N__44798\,
            I => \N__44795\
        );

    \I__9498\ : InMux
    port map (
            O => \N__44795\,
            I => \N__44791\
        );

    \I__9497\ : InMux
    port map (
            O => \N__44794\,
            I => \N__44788\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__44791\,
            I => \N__44785\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__44788\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__9494\ : Odrv12
    port map (
            O => \N__44785\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__9493\ : InMux
    port map (
            O => \N__44780\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__9492\ : CascadeMux
    port map (
            O => \N__44777\,
            I => \N__44773\
        );

    \I__9491\ : CascadeMux
    port map (
            O => \N__44776\,
            I => \N__44770\
        );

    \I__9490\ : InMux
    port map (
            O => \N__44773\,
            I => \N__44765\
        );

    \I__9489\ : InMux
    port map (
            O => \N__44770\,
            I => \N__44765\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__44765\,
            I => \N__44761\
        );

    \I__9487\ : InMux
    port map (
            O => \N__44764\,
            I => \N__44758\
        );

    \I__9486\ : Span4Mux_h
    port map (
            O => \N__44761\,
            I => \N__44755\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__44758\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__9484\ : Odrv4
    port map (
            O => \N__44755\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__9483\ : InMux
    port map (
            O => \N__44750\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__9482\ : CascadeMux
    port map (
            O => \N__44747\,
            I => \N__44743\
        );

    \I__9481\ : CascadeMux
    port map (
            O => \N__44746\,
            I => \N__44740\
        );

    \I__9480\ : InMux
    port map (
            O => \N__44743\,
            I => \N__44735\
        );

    \I__9479\ : InMux
    port map (
            O => \N__44740\,
            I => \N__44735\
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__44735\,
            I => \N__44731\
        );

    \I__9477\ : InMux
    port map (
            O => \N__44734\,
            I => \N__44728\
        );

    \I__9476\ : Span4Mux_h
    port map (
            O => \N__44731\,
            I => \N__44725\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__44728\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__9474\ : Odrv4
    port map (
            O => \N__44725\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__9473\ : InMux
    port map (
            O => \N__44720\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__9472\ : CascadeMux
    port map (
            O => \N__44717\,
            I => \N__44714\
        );

    \I__9471\ : InMux
    port map (
            O => \N__44714\,
            I => \N__44710\
        );

    \I__9470\ : InMux
    port map (
            O => \N__44713\,
            I => \N__44707\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__44710\,
            I => \N__44701\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__44707\,
            I => \N__44701\
        );

    \I__9467\ : InMux
    port map (
            O => \N__44706\,
            I => \N__44698\
        );

    \I__9466\ : Span4Mux_v
    port map (
            O => \N__44701\,
            I => \N__44695\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__44698\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__9464\ : Odrv4
    port map (
            O => \N__44695\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__9463\ : InMux
    port map (
            O => \N__44690\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__9462\ : InMux
    port map (
            O => \N__44687\,
            I => \N__44681\
        );

    \I__9461\ : InMux
    port map (
            O => \N__44686\,
            I => \N__44681\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__44681\,
            I => \N__44677\
        );

    \I__9459\ : InMux
    port map (
            O => \N__44680\,
            I => \N__44674\
        );

    \I__9458\ : Span4Mux_v
    port map (
            O => \N__44677\,
            I => \N__44671\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__44674\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__9456\ : Odrv4
    port map (
            O => \N__44671\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__9455\ : InMux
    port map (
            O => \N__44666\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__9454\ : CascadeMux
    port map (
            O => \N__44663\,
            I => \N__44660\
        );

    \I__9453\ : InMux
    port map (
            O => \N__44660\,
            I => \N__44657\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__44657\,
            I => \N__44652\
        );

    \I__9451\ : InMux
    port map (
            O => \N__44656\,
            I => \N__44649\
        );

    \I__9450\ : InMux
    port map (
            O => \N__44655\,
            I => \N__44646\
        );

    \I__9449\ : Span4Mux_h
    port map (
            O => \N__44652\,
            I => \N__44643\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__44649\,
            I => \N__44640\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__44646\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__9446\ : Odrv4
    port map (
            O => \N__44643\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__9445\ : Odrv12
    port map (
            O => \N__44640\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__9444\ : InMux
    port map (
            O => \N__44633\,
            I => \bfn_17_9_0_\
        );

    \I__9443\ : CascadeMux
    port map (
            O => \N__44630\,
            I => \N__44627\
        );

    \I__9442\ : InMux
    port map (
            O => \N__44627\,
            I => \N__44623\
        );

    \I__9441\ : CascadeMux
    port map (
            O => \N__44626\,
            I => \N__44620\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__44623\,
            I => \N__44616\
        );

    \I__9439\ : InMux
    port map (
            O => \N__44620\,
            I => \N__44613\
        );

    \I__9438\ : InMux
    port map (
            O => \N__44619\,
            I => \N__44610\
        );

    \I__9437\ : Span4Mux_h
    port map (
            O => \N__44616\,
            I => \N__44607\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__44613\,
            I => \N__44604\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__44610\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__9434\ : Odrv4
    port map (
            O => \N__44607\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__9433\ : Odrv12
    port map (
            O => \N__44604\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__9432\ : InMux
    port map (
            O => \N__44597\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__9431\ : InMux
    port map (
            O => \N__44594\,
            I => \N__44588\
        );

    \I__9430\ : InMux
    port map (
            O => \N__44593\,
            I => \N__44588\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__44588\,
            I => \N__44584\
        );

    \I__9428\ : InMux
    port map (
            O => \N__44587\,
            I => \N__44581\
        );

    \I__9427\ : Span4Mux_h
    port map (
            O => \N__44584\,
            I => \N__44578\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__44581\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__9425\ : Odrv4
    port map (
            O => \N__44578\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__9424\ : InMux
    port map (
            O => \N__44573\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__9423\ : InMux
    port map (
            O => \N__44570\,
            I => \N__44564\
        );

    \I__9422\ : InMux
    port map (
            O => \N__44569\,
            I => \N__44564\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__44564\,
            I => \N__44560\
        );

    \I__9420\ : InMux
    port map (
            O => \N__44563\,
            I => \N__44557\
        );

    \I__9419\ : Span4Mux_h
    port map (
            O => \N__44560\,
            I => \N__44554\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__44557\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__9417\ : Odrv4
    port map (
            O => \N__44554\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__9416\ : InMux
    port map (
            O => \N__44549\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__9415\ : InMux
    port map (
            O => \N__44546\,
            I => \N__44540\
        );

    \I__9414\ : InMux
    port map (
            O => \N__44545\,
            I => \N__44540\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__44540\,
            I => \N__44536\
        );

    \I__9412\ : InMux
    port map (
            O => \N__44539\,
            I => \N__44533\
        );

    \I__9411\ : Span4Mux_s2_v
    port map (
            O => \N__44536\,
            I => \N__44530\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__44533\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9409\ : Odrv4
    port map (
            O => \N__44530\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9408\ : InMux
    port map (
            O => \N__44525\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__9407\ : CascadeMux
    port map (
            O => \N__44522\,
            I => \N__44518\
        );

    \I__9406\ : CascadeMux
    port map (
            O => \N__44521\,
            I => \N__44515\
        );

    \I__9405\ : InMux
    port map (
            O => \N__44518\,
            I => \N__44510\
        );

    \I__9404\ : InMux
    port map (
            O => \N__44515\,
            I => \N__44510\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__44510\,
            I => \N__44506\
        );

    \I__9402\ : InMux
    port map (
            O => \N__44509\,
            I => \N__44503\
        );

    \I__9401\ : Span4Mux_s2_v
    port map (
            O => \N__44506\,
            I => \N__44500\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__44503\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9399\ : Odrv4
    port map (
            O => \N__44500\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9398\ : InMux
    port map (
            O => \N__44495\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__9397\ : CascadeMux
    port map (
            O => \N__44492\,
            I => \N__44488\
        );

    \I__9396\ : CascadeMux
    port map (
            O => \N__44491\,
            I => \N__44485\
        );

    \I__9395\ : InMux
    port map (
            O => \N__44488\,
            I => \N__44480\
        );

    \I__9394\ : InMux
    port map (
            O => \N__44485\,
            I => \N__44480\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__44480\,
            I => \N__44476\
        );

    \I__9392\ : InMux
    port map (
            O => \N__44479\,
            I => \N__44473\
        );

    \I__9391\ : Span4Mux_s2_v
    port map (
            O => \N__44476\,
            I => \N__44470\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__44473\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9389\ : Odrv4
    port map (
            O => \N__44470\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9388\ : InMux
    port map (
            O => \N__44465\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__9387\ : CascadeMux
    port map (
            O => \N__44462\,
            I => \N__44459\
        );

    \I__9386\ : InMux
    port map (
            O => \N__44459\,
            I => \N__44455\
        );

    \I__9385\ : InMux
    port map (
            O => \N__44458\,
            I => \N__44452\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__44455\,
            I => \N__44446\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__44452\,
            I => \N__44446\
        );

    \I__9382\ : InMux
    port map (
            O => \N__44451\,
            I => \N__44443\
        );

    \I__9381\ : Span4Mux_s3_v
    port map (
            O => \N__44446\,
            I => \N__44440\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__44443\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9379\ : Odrv4
    port map (
            O => \N__44440\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9378\ : InMux
    port map (
            O => \N__44435\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__9377\ : CascadeMux
    port map (
            O => \N__44432\,
            I => \N__44429\
        );

    \I__9376\ : InMux
    port map (
            O => \N__44429\,
            I => \N__44425\
        );

    \I__9375\ : InMux
    port map (
            O => \N__44428\,
            I => \N__44422\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__44425\,
            I => \N__44416\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__44422\,
            I => \N__44416\
        );

    \I__9372\ : InMux
    port map (
            O => \N__44421\,
            I => \N__44413\
        );

    \I__9371\ : Span4Mux_s3_v
    port map (
            O => \N__44416\,
            I => \N__44410\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__44413\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__9369\ : Odrv4
    port map (
            O => \N__44410\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__9368\ : InMux
    port map (
            O => \N__44405\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__9367\ : CascadeMux
    port map (
            O => \N__44402\,
            I => \N__44399\
        );

    \I__9366\ : InMux
    port map (
            O => \N__44399\,
            I => \N__44396\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__44396\,
            I => \N__44391\
        );

    \I__9364\ : InMux
    port map (
            O => \N__44395\,
            I => \N__44388\
        );

    \I__9363\ : InMux
    port map (
            O => \N__44394\,
            I => \N__44385\
        );

    \I__9362\ : Span4Mux_h
    port map (
            O => \N__44391\,
            I => \N__44382\
        );

    \I__9361\ : LocalMux
    port map (
            O => \N__44388\,
            I => \N__44379\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__44385\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9359\ : Odrv4
    port map (
            O => \N__44382\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9358\ : Odrv12
    port map (
            O => \N__44379\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9357\ : InMux
    port map (
            O => \N__44372\,
            I => \bfn_17_8_0_\
        );

    \I__9356\ : CascadeMux
    port map (
            O => \N__44369\,
            I => \N__44366\
        );

    \I__9355\ : InMux
    port map (
            O => \N__44366\,
            I => \N__44363\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__44363\,
            I => \N__44358\
        );

    \I__9353\ : InMux
    port map (
            O => \N__44362\,
            I => \N__44355\
        );

    \I__9352\ : InMux
    port map (
            O => \N__44361\,
            I => \N__44352\
        );

    \I__9351\ : Sp12to4
    port map (
            O => \N__44358\,
            I => \N__44347\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__44355\,
            I => \N__44347\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__44352\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__9348\ : Odrv12
    port map (
            O => \N__44347\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__9347\ : InMux
    port map (
            O => \N__44342\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__9346\ : InMux
    port map (
            O => \N__44339\,
            I => \N__44333\
        );

    \I__9345\ : InMux
    port map (
            O => \N__44338\,
            I => \N__44333\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__44333\,
            I => \N__44329\
        );

    \I__9343\ : InMux
    port map (
            O => \N__44332\,
            I => \N__44326\
        );

    \I__9342\ : Span4Mux_h
    port map (
            O => \N__44329\,
            I => \N__44323\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__44326\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__9340\ : Odrv4
    port map (
            O => \N__44323\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__9339\ : InMux
    port map (
            O => \N__44318\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__9338\ : InMux
    port map (
            O => \N__44315\,
            I => \N__44309\
        );

    \I__9337\ : InMux
    port map (
            O => \N__44314\,
            I => \N__44309\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__44309\,
            I => \N__44305\
        );

    \I__9335\ : InMux
    port map (
            O => \N__44308\,
            I => \N__44302\
        );

    \I__9334\ : Span4Mux_h
    port map (
            O => \N__44305\,
            I => \N__44299\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__44302\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__9332\ : Odrv4
    port map (
            O => \N__44299\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__9331\ : InMux
    port map (
            O => \N__44294\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__9330\ : InMux
    port map (
            O => \N__44291\,
            I => \N__44288\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__44288\,
            I => \N__44285\
        );

    \I__9328\ : Span4Mux_h
    port map (
            O => \N__44285\,
            I => \N__44281\
        );

    \I__9327\ : InMux
    port map (
            O => \N__44284\,
            I => \N__44278\
        );

    \I__9326\ : Odrv4
    port map (
            O => \N__44281\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__44278\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__9324\ : InMux
    port map (
            O => \N__44273\,
            I => \bfn_17_6_0_\
        );

    \I__9323\ : InMux
    port map (
            O => \N__44270\,
            I => \N__44267\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__44267\,
            I => \N__44264\
        );

    \I__9321\ : Span4Mux_v
    port map (
            O => \N__44264\,
            I => \N__44260\
        );

    \I__9320\ : InMux
    port map (
            O => \N__44263\,
            I => \N__44257\
        );

    \I__9319\ : Odrv4
    port map (
            O => \N__44260\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__44257\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9317\ : InMux
    port map (
            O => \N__44252\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__9316\ : InMux
    port map (
            O => \N__44249\,
            I => \N__44245\
        );

    \I__9315\ : InMux
    port map (
            O => \N__44248\,
            I => \N__44242\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__44245\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__44242\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__9312\ : InMux
    port map (
            O => \N__44237\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__9311\ : InMux
    port map (
            O => \N__44234\,
            I => \N__44231\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__44231\,
            I => \N__44227\
        );

    \I__9309\ : InMux
    port map (
            O => \N__44230\,
            I => \N__44224\
        );

    \I__9308\ : Odrv4
    port map (
            O => \N__44227\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__9307\ : LocalMux
    port map (
            O => \N__44224\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__9306\ : InMux
    port map (
            O => \N__44219\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__9305\ : InMux
    port map (
            O => \N__44216\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__9304\ : InMux
    port map (
            O => \N__44213\,
            I => \N__44210\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__44210\,
            I => \N__44206\
        );

    \I__9302\ : InMux
    port map (
            O => \N__44209\,
            I => \N__44203\
        );

    \I__9301\ : Span4Mux_h
    port map (
            O => \N__44206\,
            I => \N__44198\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__44203\,
            I => \N__44198\
        );

    \I__9299\ : Odrv4
    port map (
            O => \N__44198\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__9298\ : CEMux
    port map (
            O => \N__44195\,
            I => \N__44189\
        );

    \I__9297\ : CEMux
    port map (
            O => \N__44194\,
            I => \N__44186\
        );

    \I__9296\ : CEMux
    port map (
            O => \N__44193\,
            I => \N__44183\
        );

    \I__9295\ : CEMux
    port map (
            O => \N__44192\,
            I => \N__44179\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__44189\,
            I => \N__44176\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__44186\,
            I => \N__44171\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__44183\,
            I => \N__44171\
        );

    \I__9291\ : CEMux
    port map (
            O => \N__44182\,
            I => \N__44168\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__44179\,
            I => \N__44165\
        );

    \I__9289\ : Span4Mux_v
    port map (
            O => \N__44176\,
            I => \N__44158\
        );

    \I__9288\ : Span4Mux_v
    port map (
            O => \N__44171\,
            I => \N__44158\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__44168\,
            I => \N__44158\
        );

    \I__9286\ : Span4Mux_v
    port map (
            O => \N__44165\,
            I => \N__44153\
        );

    \I__9285\ : Span4Mux_h
    port map (
            O => \N__44158\,
            I => \N__44153\
        );

    \I__9284\ : Odrv4
    port map (
            O => \N__44153\,
            I => \delay_measurement_inst.delay_hc_timer.N_165_i\
        );

    \I__9283\ : InMux
    port map (
            O => \N__44150\,
            I => \N__44146\
        );

    \I__9282\ : InMux
    port map (
            O => \N__44149\,
            I => \N__44143\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__44146\,
            I => \N__44139\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__44143\,
            I => \N__44136\
        );

    \I__9279\ : InMux
    port map (
            O => \N__44142\,
            I => \N__44133\
        );

    \I__9278\ : Odrv4
    port map (
            O => \N__44139\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9277\ : Odrv12
    port map (
            O => \N__44136\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__44133\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9275\ : InMux
    port map (
            O => \N__44126\,
            I => \bfn_17_7_0_\
        );

    \I__9274\ : CascadeMux
    port map (
            O => \N__44123\,
            I => \N__44120\
        );

    \I__9273\ : InMux
    port map (
            O => \N__44120\,
            I => \N__44116\
        );

    \I__9272\ : InMux
    port map (
            O => \N__44119\,
            I => \N__44112\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__44116\,
            I => \N__44109\
        );

    \I__9270\ : InMux
    port map (
            O => \N__44115\,
            I => \N__44106\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__44112\,
            I => \N__44101\
        );

    \I__9268\ : Span4Mux_s2_v
    port map (
            O => \N__44109\,
            I => \N__44101\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__44106\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__9266\ : Odrv4
    port map (
            O => \N__44101\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__9265\ : InMux
    port map (
            O => \N__44096\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__9264\ : CascadeMux
    port map (
            O => \N__44093\,
            I => \N__44089\
        );

    \I__9263\ : InMux
    port map (
            O => \N__44092\,
            I => \N__44086\
        );

    \I__9262\ : InMux
    port map (
            O => \N__44089\,
            I => \N__44083\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__44086\,
            I => \N__44077\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__44083\,
            I => \N__44077\
        );

    \I__9259\ : InMux
    port map (
            O => \N__44082\,
            I => \N__44074\
        );

    \I__9258\ : Span4Mux_s2_v
    port map (
            O => \N__44077\,
            I => \N__44071\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__44074\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9256\ : Odrv4
    port map (
            O => \N__44071\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9255\ : InMux
    port map (
            O => \N__44066\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__9254\ : InMux
    port map (
            O => \N__44063\,
            I => \N__44060\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__44060\,
            I => \N__44057\
        );

    \I__9252\ : Span4Mux_h
    port map (
            O => \N__44057\,
            I => \N__44053\
        );

    \I__9251\ : InMux
    port map (
            O => \N__44056\,
            I => \N__44050\
        );

    \I__9250\ : Odrv4
    port map (
            O => \N__44053\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__44050\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__9248\ : InMux
    port map (
            O => \N__44045\,
            I => \bfn_17_5_0_\
        );

    \I__9247\ : InMux
    port map (
            O => \N__44042\,
            I => \N__44039\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__44039\,
            I => \N__44036\
        );

    \I__9245\ : Span4Mux_h
    port map (
            O => \N__44036\,
            I => \N__44032\
        );

    \I__9244\ : InMux
    port map (
            O => \N__44035\,
            I => \N__44029\
        );

    \I__9243\ : Odrv4
    port map (
            O => \N__44032\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__44029\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9241\ : InMux
    port map (
            O => \N__44024\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__9240\ : InMux
    port map (
            O => \N__44021\,
            I => \N__44018\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__44018\,
            I => \N__44015\
        );

    \I__9238\ : Span4Mux_v
    port map (
            O => \N__44015\,
            I => \N__44011\
        );

    \I__9237\ : InMux
    port map (
            O => \N__44014\,
            I => \N__44008\
        );

    \I__9236\ : Odrv4
    port map (
            O => \N__44011\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__44008\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__9234\ : InMux
    port map (
            O => \N__44003\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__9233\ : InMux
    port map (
            O => \N__44000\,
            I => \N__43996\
        );

    \I__9232\ : CascadeMux
    port map (
            O => \N__43999\,
            I => \N__43993\
        );

    \I__9231\ : LocalMux
    port map (
            O => \N__43996\,
            I => \N__43990\
        );

    \I__9230\ : InMux
    port map (
            O => \N__43993\,
            I => \N__43987\
        );

    \I__9229\ : Odrv4
    port map (
            O => \N__43990\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__43987\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9227\ : InMux
    port map (
            O => \N__43982\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__9226\ : InMux
    port map (
            O => \N__43979\,
            I => \N__43976\
        );

    \I__9225\ : LocalMux
    port map (
            O => \N__43976\,
            I => \N__43972\
        );

    \I__9224\ : CascadeMux
    port map (
            O => \N__43975\,
            I => \N__43969\
        );

    \I__9223\ : Span4Mux_h
    port map (
            O => \N__43972\,
            I => \N__43966\
        );

    \I__9222\ : InMux
    port map (
            O => \N__43969\,
            I => \N__43963\
        );

    \I__9221\ : Odrv4
    port map (
            O => \N__43966\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__43963\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9219\ : InMux
    port map (
            O => \N__43958\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__9218\ : InMux
    port map (
            O => \N__43955\,
            I => \N__43952\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__43952\,
            I => \N__43949\
        );

    \I__9216\ : Span4Mux_h
    port map (
            O => \N__43949\,
            I => \N__43945\
        );

    \I__9215\ : InMux
    port map (
            O => \N__43948\,
            I => \N__43942\
        );

    \I__9214\ : Odrv4
    port map (
            O => \N__43945\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__43942\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__9212\ : InMux
    port map (
            O => \N__43937\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__9211\ : InMux
    port map (
            O => \N__43934\,
            I => \N__43931\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__43931\,
            I => \N__43927\
        );

    \I__9209\ : CascadeMux
    port map (
            O => \N__43930\,
            I => \N__43924\
        );

    \I__9208\ : Span4Mux_v
    port map (
            O => \N__43927\,
            I => \N__43921\
        );

    \I__9207\ : InMux
    port map (
            O => \N__43924\,
            I => \N__43918\
        );

    \I__9206\ : Odrv4
    port map (
            O => \N__43921\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__43918\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__9204\ : InMux
    port map (
            O => \N__43913\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__9203\ : InMux
    port map (
            O => \N__43910\,
            I => \N__43907\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__43907\,
            I => \N__43904\
        );

    \I__9201\ : Span4Mux_h
    port map (
            O => \N__43904\,
            I => \N__43900\
        );

    \I__9200\ : InMux
    port map (
            O => \N__43903\,
            I => \N__43897\
        );

    \I__9199\ : Odrv4
    port map (
            O => \N__43900\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__43897\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__9197\ : InMux
    port map (
            O => \N__43892\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__9196\ : InMux
    port map (
            O => \N__43889\,
            I => \N__43886\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__43886\,
            I => \N__43882\
        );

    \I__9194\ : InMux
    port map (
            O => \N__43885\,
            I => \N__43879\
        );

    \I__9193\ : Span4Mux_h
    port map (
            O => \N__43882\,
            I => \N__43876\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__43879\,
            I => \N__43873\
        );

    \I__9191\ : Odrv4
    port map (
            O => \N__43876\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__9190\ : Odrv4
    port map (
            O => \N__43873\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__9189\ : InMux
    port map (
            O => \N__43868\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__9188\ : InMux
    port map (
            O => \N__43865\,
            I => \N__43862\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__43862\,
            I => \N__43859\
        );

    \I__9186\ : Span4Mux_h
    port map (
            O => \N__43859\,
            I => \N__43855\
        );

    \I__9185\ : InMux
    port map (
            O => \N__43858\,
            I => \N__43852\
        );

    \I__9184\ : Odrv4
    port map (
            O => \N__43855\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__9183\ : LocalMux
    port map (
            O => \N__43852\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__9182\ : InMux
    port map (
            O => \N__43847\,
            I => \bfn_17_4_0_\
        );

    \I__9181\ : InMux
    port map (
            O => \N__43844\,
            I => \N__43841\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__43841\,
            I => \N__43838\
        );

    \I__9179\ : Span4Mux_v
    port map (
            O => \N__43838\,
            I => \N__43834\
        );

    \I__9178\ : InMux
    port map (
            O => \N__43837\,
            I => \N__43831\
        );

    \I__9177\ : Odrv4
    port map (
            O => \N__43834\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__43831\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__9175\ : InMux
    port map (
            O => \N__43826\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__9174\ : InMux
    port map (
            O => \N__43823\,
            I => \N__43820\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__43820\,
            I => \N__43817\
        );

    \I__9172\ : Span4Mux_h
    port map (
            O => \N__43817\,
            I => \N__43813\
        );

    \I__9171\ : InMux
    port map (
            O => \N__43816\,
            I => \N__43810\
        );

    \I__9170\ : Odrv4
    port map (
            O => \N__43813\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__43810\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__9168\ : InMux
    port map (
            O => \N__43805\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__9167\ : InMux
    port map (
            O => \N__43802\,
            I => \N__43799\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__43799\,
            I => \N__43796\
        );

    \I__9165\ : Span4Mux_h
    port map (
            O => \N__43796\,
            I => \N__43792\
        );

    \I__9164\ : InMux
    port map (
            O => \N__43795\,
            I => \N__43789\
        );

    \I__9163\ : Odrv4
    port map (
            O => \N__43792\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__43789\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__9161\ : InMux
    port map (
            O => \N__43784\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__9160\ : InMux
    port map (
            O => \N__43781\,
            I => \N__43778\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__43778\,
            I => \N__43775\
        );

    \I__9158\ : Span4Mux_h
    port map (
            O => \N__43775\,
            I => \N__43771\
        );

    \I__9157\ : InMux
    port map (
            O => \N__43774\,
            I => \N__43768\
        );

    \I__9156\ : Odrv4
    port map (
            O => \N__43771\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__43768\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__9154\ : InMux
    port map (
            O => \N__43763\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__9153\ : InMux
    port map (
            O => \N__43760\,
            I => \N__43757\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__43757\,
            I => \N__43753\
        );

    \I__9151\ : InMux
    port map (
            O => \N__43756\,
            I => \N__43750\
        );

    \I__9150\ : Odrv4
    port map (
            O => \N__43753\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__43750\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__9148\ : InMux
    port map (
            O => \N__43745\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__9147\ : InMux
    port map (
            O => \N__43742\,
            I => \N__43739\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__43739\,
            I => \N__43736\
        );

    \I__9145\ : Span4Mux_v
    port map (
            O => \N__43736\,
            I => \N__43733\
        );

    \I__9144\ : Span4Mux_h
    port map (
            O => \N__43733\,
            I => \N__43729\
        );

    \I__9143\ : InMux
    port map (
            O => \N__43732\,
            I => \N__43726\
        );

    \I__9142\ : Odrv4
    port map (
            O => \N__43729\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__43726\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__9140\ : InMux
    port map (
            O => \N__43721\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__9139\ : InMux
    port map (
            O => \N__43718\,
            I => \N__43715\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__43715\,
            I => \N__43711\
        );

    \I__9137\ : CascadeMux
    port map (
            O => \N__43714\,
            I => \N__43708\
        );

    \I__9136\ : Span4Mux_v
    port map (
            O => \N__43711\,
            I => \N__43705\
        );

    \I__9135\ : InMux
    port map (
            O => \N__43708\,
            I => \N__43702\
        );

    \I__9134\ : Odrv4
    port map (
            O => \N__43705\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__43702\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__9132\ : InMux
    port map (
            O => \N__43697\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__9131\ : InMux
    port map (
            O => \N__43694\,
            I => \N__43691\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__43691\,
            I => \N__43688\
        );

    \I__9129\ : Span4Mux_v
    port map (
            O => \N__43688\,
            I => \N__43684\
        );

    \I__9128\ : InMux
    port map (
            O => \N__43687\,
            I => \N__43681\
        );

    \I__9127\ : Odrv4
    port map (
            O => \N__43684\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__43681\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__9125\ : InMux
    port map (
            O => \N__43676\,
            I => \N__43673\
        );

    \I__9124\ : LocalMux
    port map (
            O => \N__43673\,
            I => \N__43670\
        );

    \I__9123\ : Span4Mux_v
    port map (
            O => \N__43670\,
            I => \N__43666\
        );

    \I__9122\ : InMux
    port map (
            O => \N__43669\,
            I => \N__43663\
        );

    \I__9121\ : Odrv4
    port map (
            O => \N__43666\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__43663\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__9119\ : InMux
    port map (
            O => \N__43658\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__9118\ : InMux
    port map (
            O => \N__43655\,
            I => \N__43652\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__43652\,
            I => \N__43649\
        );

    \I__9116\ : Span4Mux_h
    port map (
            O => \N__43649\,
            I => \N__43645\
        );

    \I__9115\ : InMux
    port map (
            O => \N__43648\,
            I => \N__43642\
        );

    \I__9114\ : Odrv4
    port map (
            O => \N__43645\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__43642\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__9112\ : InMux
    port map (
            O => \N__43637\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__9111\ : InMux
    port map (
            O => \N__43634\,
            I => \N__43631\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__43631\,
            I => \N__43628\
        );

    \I__9109\ : Span4Mux_h
    port map (
            O => \N__43628\,
            I => \N__43624\
        );

    \I__9108\ : InMux
    port map (
            O => \N__43627\,
            I => \N__43621\
        );

    \I__9107\ : Odrv4
    port map (
            O => \N__43624\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__43621\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__9105\ : InMux
    port map (
            O => \N__43616\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__9104\ : CascadeMux
    port map (
            O => \N__43613\,
            I => \N__43609\
        );

    \I__9103\ : InMux
    port map (
            O => \N__43612\,
            I => \N__43606\
        );

    \I__9102\ : InMux
    port map (
            O => \N__43609\,
            I => \N__43603\
        );

    \I__9101\ : LocalMux
    port map (
            O => \N__43606\,
            I => \N__43600\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__43603\,
            I => \N__43597\
        );

    \I__9099\ : Span4Mux_h
    port map (
            O => \N__43600\,
            I => \N__43594\
        );

    \I__9098\ : Span4Mux_h
    port map (
            O => \N__43597\,
            I => \N__43591\
        );

    \I__9097\ : Odrv4
    port map (
            O => \N__43594\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__9096\ : Odrv4
    port map (
            O => \N__43591\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__9095\ : InMux
    port map (
            O => \N__43586\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__9094\ : InMux
    port map (
            O => \N__43583\,
            I => \N__43579\
        );

    \I__9093\ : InMux
    port map (
            O => \N__43582\,
            I => \N__43576\
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__43579\,
            I => \N__43573\
        );

    \I__9091\ : LocalMux
    port map (
            O => \N__43576\,
            I => \N__43570\
        );

    \I__9090\ : Span4Mux_h
    port map (
            O => \N__43573\,
            I => \N__43567\
        );

    \I__9089\ : Span4Mux_h
    port map (
            O => \N__43570\,
            I => \N__43564\
        );

    \I__9088\ : Odrv4
    port map (
            O => \N__43567\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__9087\ : Odrv4
    port map (
            O => \N__43564\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__9086\ : InMux
    port map (
            O => \N__43559\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__9085\ : InMux
    port map (
            O => \N__43556\,
            I => \N__43553\
        );

    \I__9084\ : LocalMux
    port map (
            O => \N__43553\,
            I => \N__43549\
        );

    \I__9083\ : CascadeMux
    port map (
            O => \N__43552\,
            I => \N__43546\
        );

    \I__9082\ : Span4Mux_v
    port map (
            O => \N__43549\,
            I => \N__43543\
        );

    \I__9081\ : InMux
    port map (
            O => \N__43546\,
            I => \N__43540\
        );

    \I__9080\ : Span4Mux_h
    port map (
            O => \N__43543\,
            I => \N__43537\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__43540\,
            I => \N__43534\
        );

    \I__9078\ : Odrv4
    port map (
            O => \N__43537\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__9077\ : Odrv4
    port map (
            O => \N__43534\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__9076\ : InMux
    port map (
            O => \N__43529\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__9075\ : InMux
    port map (
            O => \N__43526\,
            I => \N__43523\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__43523\,
            I => \N__43520\
        );

    \I__9073\ : Span4Mux_s1_h
    port map (
            O => \N__43520\,
            I => \N__43516\
        );

    \I__9072\ : InMux
    port map (
            O => \N__43519\,
            I => \N__43513\
        );

    \I__9071\ : Span4Mux_h
    port map (
            O => \N__43516\,
            I => \N__43510\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__43513\,
            I => \N__43505\
        );

    \I__9069\ : Span4Mux_h
    port map (
            O => \N__43510\,
            I => \N__43505\
        );

    \I__9068\ : Odrv4
    port map (
            O => \N__43505\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__9067\ : InMux
    port map (
            O => \N__43502\,
            I => \N__43499\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__43499\,
            I => \N__43496\
        );

    \I__9065\ : Sp12to4
    port map (
            O => \N__43496\,
            I => \N__43492\
        );

    \I__9064\ : InMux
    port map (
            O => \N__43495\,
            I => \N__43489\
        );

    \I__9063\ : Span12Mux_v
    port map (
            O => \N__43492\,
            I => \N__43486\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__43489\,
            I => \N__43483\
        );

    \I__9061\ : Span12Mux_h
    port map (
            O => \N__43486\,
            I => \N__43480\
        );

    \I__9060\ : Odrv4
    port map (
            O => \N__43483\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__9059\ : Odrv12
    port map (
            O => \N__43480\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__9058\ : InMux
    port map (
            O => \N__43475\,
            I => \N__43472\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__43472\,
            I => \N__43469\
        );

    \I__9056\ : Span4Mux_v
    port map (
            O => \N__43469\,
            I => \N__43466\
        );

    \I__9055\ : Span4Mux_v
    port map (
            O => \N__43466\,
            I => \N__43463\
        );

    \I__9054\ : Span4Mux_v
    port map (
            O => \N__43463\,
            I => \N__43459\
        );

    \I__9053\ : InMux
    port map (
            O => \N__43462\,
            I => \N__43456\
        );

    \I__9052\ : Sp12to4
    port map (
            O => \N__43459\,
            I => \N__43453\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__43456\,
            I => \N__43450\
        );

    \I__9050\ : Span12Mux_s9_h
    port map (
            O => \N__43453\,
            I => \N__43447\
        );

    \I__9049\ : Odrv4
    port map (
            O => \N__43450\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__9048\ : Odrv12
    port map (
            O => \N__43447\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__9047\ : InMux
    port map (
            O => \N__43442\,
            I => \N__43439\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__43439\,
            I => \N__43436\
        );

    \I__9045\ : Span12Mux_v
    port map (
            O => \N__43436\,
            I => \N__43432\
        );

    \I__9044\ : InMux
    port map (
            O => \N__43435\,
            I => \N__43429\
        );

    \I__9043\ : Span12Mux_h
    port map (
            O => \N__43432\,
            I => \N__43426\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__43429\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__9041\ : Odrv12
    port map (
            O => \N__43426\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__9040\ : InMux
    port map (
            O => \N__43421\,
            I => \N__43418\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__43418\,
            I => \N__43415\
        );

    \I__9038\ : Span4Mux_s2_h
    port map (
            O => \N__43415\,
            I => \N__43412\
        );

    \I__9037\ : Span4Mux_h
    port map (
            O => \N__43412\,
            I => \N__43408\
        );

    \I__9036\ : InMux
    port map (
            O => \N__43411\,
            I => \N__43405\
        );

    \I__9035\ : Span4Mux_v
    port map (
            O => \N__43408\,
            I => \N__43402\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__43405\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__9033\ : Odrv4
    port map (
            O => \N__43402\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__9032\ : InMux
    port map (
            O => \N__43397\,
            I => \N__43394\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__43394\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\
        );

    \I__9030\ : InMux
    port map (
            O => \N__43391\,
            I => \N__43388\
        );

    \I__9029\ : LocalMux
    port map (
            O => \N__43388\,
            I => \N__43385\
        );

    \I__9028\ : Span4Mux_s2_h
    port map (
            O => \N__43385\,
            I => \N__43382\
        );

    \I__9027\ : Sp12to4
    port map (
            O => \N__43382\,
            I => \N__43378\
        );

    \I__9026\ : InMux
    port map (
            O => \N__43381\,
            I => \N__43375\
        );

    \I__9025\ : Span12Mux_h
    port map (
            O => \N__43378\,
            I => \N__43372\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__43375\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__9023\ : Odrv12
    port map (
            O => \N__43372\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__9022\ : InMux
    port map (
            O => \N__43367\,
            I => \N__43364\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__43364\,
            I => \N__43361\
        );

    \I__9020\ : Span12Mux_s7_h
    port map (
            O => \N__43361\,
            I => \N__43357\
        );

    \I__9019\ : InMux
    port map (
            O => \N__43360\,
            I => \N__43354\
        );

    \I__9018\ : Span12Mux_v
    port map (
            O => \N__43357\,
            I => \N__43351\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__43354\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__9016\ : Odrv12
    port map (
            O => \N__43351\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__9015\ : InMux
    port map (
            O => \N__43346\,
            I => \N__43343\
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__43343\,
            I => \N__43340\
        );

    \I__9013\ : Span12Mux_v
    port map (
            O => \N__43340\,
            I => \N__43336\
        );

    \I__9012\ : InMux
    port map (
            O => \N__43339\,
            I => \N__43333\
        );

    \I__9011\ : Span12Mux_h
    port map (
            O => \N__43336\,
            I => \N__43330\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__43333\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__9009\ : Odrv12
    port map (
            O => \N__43330\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__9008\ : InMux
    port map (
            O => \N__43325\,
            I => \N__43322\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__43322\,
            I => \N__43319\
        );

    \I__9006\ : Span4Mux_v
    port map (
            O => \N__43319\,
            I => \N__43316\
        );

    \I__9005\ : Span4Mux_v
    port map (
            O => \N__43316\,
            I => \N__43313\
        );

    \I__9004\ : Sp12to4
    port map (
            O => \N__43313\,
            I => \N__43310\
        );

    \I__9003\ : Span12Mux_s3_h
    port map (
            O => \N__43310\,
            I => \N__43306\
        );

    \I__9002\ : InMux
    port map (
            O => \N__43309\,
            I => \N__43303\
        );

    \I__9001\ : Span12Mux_h
    port map (
            O => \N__43306\,
            I => \N__43300\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__43303\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__8999\ : Odrv12
    port map (
            O => \N__43300\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__8998\ : InMux
    port map (
            O => \N__43295\,
            I => \N__43292\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__43292\,
            I => \N__43289\
        );

    \I__8996\ : Span4Mux_v
    port map (
            O => \N__43289\,
            I => \N__43286\
        );

    \I__8995\ : Odrv4
    port map (
            O => \N__43286\,
            I => \current_shift_inst.un38_control_input_0_s1_13\
        );

    \I__8994\ : InMux
    port map (
            O => \N__43283\,
            I => \N__43280\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__43280\,
            I => \N__43277\
        );

    \I__8992\ : Odrv12
    port map (
            O => \N__43277\,
            I => \current_shift_inst.un38_control_input_0_s1_14\
        );

    \I__8991\ : InMux
    port map (
            O => \N__43274\,
            I => \N__43271\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__43271\,
            I => \N__43268\
        );

    \I__8989\ : Span4Mux_v
    port map (
            O => \N__43268\,
            I => \N__43265\
        );

    \I__8988\ : Odrv4
    port map (
            O => \N__43265\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__8987\ : InMux
    port map (
            O => \N__43262\,
            I => \N__43259\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__43259\,
            I => \N__43256\
        );

    \I__8985\ : Odrv12
    port map (
            O => \N__43256\,
            I => \current_shift_inst.un38_control_input_0_s1_11\
        );

    \I__8984\ : InMux
    port map (
            O => \N__43253\,
            I => \N__43250\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__43250\,
            I => \N__43247\
        );

    \I__8982\ : Odrv12
    port map (
            O => \N__43247\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__8981\ : InMux
    port map (
            O => \N__43244\,
            I => \N__43241\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__43241\,
            I => \N__43238\
        );

    \I__8979\ : Odrv12
    port map (
            O => \N__43238\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__8978\ : InMux
    port map (
            O => \N__43235\,
            I => \N__43232\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__43232\,
            I => \N__43229\
        );

    \I__8976\ : Span4Mux_v
    port map (
            O => \N__43229\,
            I => \N__43226\
        );

    \I__8975\ : Odrv4
    port map (
            O => \N__43226\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__8974\ : InMux
    port map (
            O => \N__43223\,
            I => \N__43220\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__43220\,
            I => \N__43217\
        );

    \I__8972\ : Span4Mux_v
    port map (
            O => \N__43217\,
            I => \N__43214\
        );

    \I__8971\ : Odrv4
    port map (
            O => \N__43214\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__8970\ : CascadeMux
    port map (
            O => \N__43211\,
            I => \N__43208\
        );

    \I__8969\ : InMux
    port map (
            O => \N__43208\,
            I => \N__43205\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__43205\,
            I => \N__43202\
        );

    \I__8967\ : Odrv12
    port map (
            O => \N__43202\,
            I => \current_shift_inst.un38_control_input_0_s1_18\
        );

    \I__8966\ : InMux
    port map (
            O => \N__43199\,
            I => \N__43196\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__43196\,
            I => \N__43193\
        );

    \I__8964\ : Span4Mux_v
    port map (
            O => \N__43193\,
            I => \N__43190\
        );

    \I__8963\ : Odrv4
    port map (
            O => \N__43190\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__8962\ : InMux
    port map (
            O => \N__43187\,
            I => \N__43184\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__43184\,
            I => \N__43181\
        );

    \I__8960\ : Odrv12
    port map (
            O => \N__43181\,
            I => \current_shift_inst.un38_control_input_0_s1_7\
        );

    \I__8959\ : InMux
    port map (
            O => \N__43178\,
            I => \N__43175\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__43175\,
            I => \N__43172\
        );

    \I__8957\ : Span12Mux_v
    port map (
            O => \N__43172\,
            I => \N__43169\
        );

    \I__8956\ : Odrv12
    port map (
            O => \N__43169\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__8955\ : InMux
    port map (
            O => \N__43166\,
            I => \N__43163\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__43163\,
            I => \N__43160\
        );

    \I__8953\ : Odrv12
    port map (
            O => \N__43160\,
            I => \current_shift_inst.un38_control_input_0_s1_10\
        );

    \I__8952\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43154\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__43154\,
            I => \N__43151\
        );

    \I__8950\ : Odrv12
    port map (
            O => \N__43151\,
            I => \current_shift_inst.un38_control_input_0_s1_9\
        );

    \I__8949\ : InMux
    port map (
            O => \N__43148\,
            I => \N__43145\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__43145\,
            I => \N__43142\
        );

    \I__8947\ : Odrv12
    port map (
            O => \N__43142\,
            I => \current_shift_inst.un38_control_input_0_s1_8\
        );

    \I__8946\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43136\
        );

    \I__8945\ : LocalMux
    port map (
            O => \N__43136\,
            I => \N__43133\
        );

    \I__8944\ : Span4Mux_v
    port map (
            O => \N__43133\,
            I => \N__43130\
        );

    \I__8943\ : Odrv4
    port map (
            O => \N__43130\,
            I => \current_shift_inst.un38_control_input_0_s1_12\
        );

    \I__8942\ : InMux
    port map (
            O => \N__43127\,
            I => \N__43124\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__43124\,
            I => \N__43121\
        );

    \I__8940\ : Odrv12
    port map (
            O => \N__43121\,
            I => \current_shift_inst.un38_control_input_0_s1_3\
        );

    \I__8939\ : CascadeMux
    port map (
            O => \N__43118\,
            I => \current_shift_inst.control_input_axb_0_cascade_\
        );

    \I__8938\ : CascadeMux
    port map (
            O => \N__43115\,
            I => \N__43112\
        );

    \I__8937\ : InMux
    port map (
            O => \N__43112\,
            I => \N__43109\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__43109\,
            I => \N__43104\
        );

    \I__8935\ : InMux
    port map (
            O => \N__43108\,
            I => \N__43101\
        );

    \I__8934\ : InMux
    port map (
            O => \N__43107\,
            I => \N__43098\
        );

    \I__8933\ : Span4Mux_v
    port map (
            O => \N__43104\,
            I => \N__43095\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__43101\,
            I => \N__43092\
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__43098\,
            I => \N__43089\
        );

    \I__8930\ : Span4Mux_v
    port map (
            O => \N__43095\,
            I => \N__43085\
        );

    \I__8929\ : Sp12to4
    port map (
            O => \N__43092\,
            I => \N__43082\
        );

    \I__8928\ : Span4Mux_v
    port map (
            O => \N__43089\,
            I => \N__43079\
        );

    \I__8927\ : InMux
    port map (
            O => \N__43088\,
            I => \N__43076\
        );

    \I__8926\ : Odrv4
    port map (
            O => \N__43085\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8925\ : Odrv12
    port map (
            O => \N__43082\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8924\ : Odrv4
    port map (
            O => \N__43079\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__43076\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8922\ : InMux
    port map (
            O => \N__43067\,
            I => \N__43063\
        );

    \I__8921\ : CascadeMux
    port map (
            O => \N__43066\,
            I => \N__43060\
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__43063\,
            I => \N__43056\
        );

    \I__8919\ : InMux
    port map (
            O => \N__43060\,
            I => \N__43053\
        );

    \I__8918\ : InMux
    port map (
            O => \N__43059\,
            I => \N__43050\
        );

    \I__8917\ : Span4Mux_v
    port map (
            O => \N__43056\,
            I => \N__43047\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__43053\,
            I => \N__43044\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__43050\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__8914\ : Odrv4
    port map (
            O => \N__43047\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__8913\ : Odrv4
    port map (
            O => \N__43044\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__8912\ : InMux
    port map (
            O => \N__43037\,
            I => \N__43034\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__43034\,
            I => \N__43031\
        );

    \I__8910\ : Odrv4
    port map (
            O => \N__43031\,
            I => \current_shift_inst.un38_control_input_0_s1_19\
        );

    \I__8909\ : InMux
    port map (
            O => \N__43028\,
            I => \N__43025\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__43025\,
            I => \N__43022\
        );

    \I__8907\ : Span12Mux_v
    port map (
            O => \N__43022\,
            I => \N__43019\
        );

    \I__8906\ : Odrv12
    port map (
            O => \N__43019\,
            I => \current_shift_inst.un38_control_input_0_s1_17\
        );

    \I__8905\ : InMux
    port map (
            O => \N__43016\,
            I => \N__43013\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__43013\,
            I => \N__43010\
        );

    \I__8903\ : Odrv12
    port map (
            O => \N__43010\,
            I => \current_shift_inst.un38_control_input_0_s1_15\
        );

    \I__8902\ : CascadeMux
    port map (
            O => \N__43007\,
            I => \N__43004\
        );

    \I__8901\ : InMux
    port map (
            O => \N__43004\,
            I => \N__43001\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__43001\,
            I => \N__42998\
        );

    \I__8899\ : Span4Mux_v
    port map (
            O => \N__42998\,
            I => \N__42995\
        );

    \I__8898\ : Odrv4
    port map (
            O => \N__42995\,
            I => \current_shift_inst.un38_control_input_0_s1_16\
        );

    \I__8897\ : CascadeMux
    port map (
            O => \N__42992\,
            I => \N__42988\
        );

    \I__8896\ : InMux
    port map (
            O => \N__42991\,
            I => \N__42984\
        );

    \I__8895\ : InMux
    port map (
            O => \N__42988\,
            I => \N__42981\
        );

    \I__8894\ : InMux
    port map (
            O => \N__42987\,
            I => \N__42978\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__42984\,
            I => \N__42975\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__42981\,
            I => \N__42972\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__42978\,
            I => \N__42969\
        );

    \I__8890\ : Span4Mux_v
    port map (
            O => \N__42975\,
            I => \N__42965\
        );

    \I__8889\ : Span4Mux_v
    port map (
            O => \N__42972\,
            I => \N__42962\
        );

    \I__8888\ : Span4Mux_v
    port map (
            O => \N__42969\,
            I => \N__42959\
        );

    \I__8887\ : InMux
    port map (
            O => \N__42968\,
            I => \N__42956\
        );

    \I__8886\ : Odrv4
    port map (
            O => \N__42965\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8885\ : Odrv4
    port map (
            O => \N__42962\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8884\ : Odrv4
    port map (
            O => \N__42959\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__42956\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8882\ : InMux
    port map (
            O => \N__42947\,
            I => \N__42944\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__42944\,
            I => \N__42939\
        );

    \I__8880\ : InMux
    port map (
            O => \N__42943\,
            I => \N__42936\
        );

    \I__8879\ : InMux
    port map (
            O => \N__42942\,
            I => \N__42933\
        );

    \I__8878\ : Span4Mux_h
    port map (
            O => \N__42939\,
            I => \N__42930\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__42936\,
            I => \N__42927\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__42933\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__8875\ : Odrv4
    port map (
            O => \N__42930\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__8874\ : Odrv12
    port map (
            O => \N__42927\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__8873\ : InMux
    port map (
            O => \N__42920\,
            I => \N__42917\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__42917\,
            I => \N__42914\
        );

    \I__8871\ : Span4Mux_v
    port map (
            O => \N__42914\,
            I => \N__42911\
        );

    \I__8870\ : Odrv4
    port map (
            O => \N__42911\,
            I => \current_shift_inst.un38_control_input_0_s1_4\
        );

    \I__8869\ : InMux
    port map (
            O => \N__42908\,
            I => \N__42905\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__42905\,
            I => \N__42902\
        );

    \I__8867\ : Span4Mux_v
    port map (
            O => \N__42902\,
            I => \N__42899\
        );

    \I__8866\ : Odrv4
    port map (
            O => \N__42899\,
            I => \current_shift_inst.un38_control_input_0_s1_5\
        );

    \I__8865\ : InMux
    port map (
            O => \N__42896\,
            I => \N__42893\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__42893\,
            I => \N__42890\
        );

    \I__8863\ : Odrv12
    port map (
            O => \N__42890\,
            I => \current_shift_inst.un38_control_input_0_s1_6\
        );

    \I__8862\ : CascadeMux
    port map (
            O => \N__42887\,
            I => \N__42884\
        );

    \I__8861\ : InMux
    port map (
            O => \N__42884\,
            I => \N__42881\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__42881\,
            I => \N__42877\
        );

    \I__8859\ : CascadeMux
    port map (
            O => \N__42880\,
            I => \N__42873\
        );

    \I__8858\ : Span4Mux_v
    port map (
            O => \N__42877\,
            I => \N__42870\
        );

    \I__8857\ : InMux
    port map (
            O => \N__42876\,
            I => \N__42867\
        );

    \I__8856\ : InMux
    port map (
            O => \N__42873\,
            I => \N__42864\
        );

    \I__8855\ : Span4Mux_h
    port map (
            O => \N__42870\,
            I => \N__42861\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__42867\,
            I => \N__42858\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__42864\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__8852\ : Odrv4
    port map (
            O => \N__42861\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__8851\ : Odrv12
    port map (
            O => \N__42858\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__8850\ : InMux
    port map (
            O => \N__42851\,
            I => \N__42847\
        );

    \I__8849\ : CascadeMux
    port map (
            O => \N__42850\,
            I => \N__42844\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__42847\,
            I => \N__42840\
        );

    \I__8847\ : InMux
    port map (
            O => \N__42844\,
            I => \N__42837\
        );

    \I__8846\ : InMux
    port map (
            O => \N__42843\,
            I => \N__42834\
        );

    \I__8845\ : Span4Mux_h
    port map (
            O => \N__42840\,
            I => \N__42829\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__42837\,
            I => \N__42829\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__42834\,
            I => \N__42825\
        );

    \I__8842\ : Span4Mux_v
    port map (
            O => \N__42829\,
            I => \N__42822\
        );

    \I__8841\ : InMux
    port map (
            O => \N__42828\,
            I => \N__42819\
        );

    \I__8840\ : Odrv12
    port map (
            O => \N__42825\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__8839\ : Odrv4
    port map (
            O => \N__42822\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__42819\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__8837\ : CascadeMux
    port map (
            O => \N__42812\,
            I => \N__42809\
        );

    \I__8836\ : InMux
    port map (
            O => \N__42809\,
            I => \N__42806\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__42806\,
            I => \N__42803\
        );

    \I__8834\ : Odrv4
    port map (
            O => \N__42803\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\
        );

    \I__8833\ : InMux
    port map (
            O => \N__42800\,
            I => \N__42797\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__42797\,
            I => \N__42793\
        );

    \I__8831\ : InMux
    port map (
            O => \N__42796\,
            I => \N__42790\
        );

    \I__8830\ : Span4Mux_v
    port map (
            O => \N__42793\,
            I => \N__42787\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__42790\,
            I => \N__42784\
        );

    \I__8828\ : Odrv4
    port map (
            O => \N__42787\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__8827\ : Odrv12
    port map (
            O => \N__42784\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__8826\ : InMux
    port map (
            O => \N__42779\,
            I => \N__42758\
        );

    \I__8825\ : CascadeMux
    port map (
            O => \N__42778\,
            I => \N__42755\
        );

    \I__8824\ : CascadeMux
    port map (
            O => \N__42777\,
            I => \N__42752\
        );

    \I__8823\ : CascadeMux
    port map (
            O => \N__42776\,
            I => \N__42749\
        );

    \I__8822\ : CascadeMux
    port map (
            O => \N__42775\,
            I => \N__42746\
        );

    \I__8821\ : CascadeMux
    port map (
            O => \N__42774\,
            I => \N__42743\
        );

    \I__8820\ : CascadeMux
    port map (
            O => \N__42773\,
            I => \N__42740\
        );

    \I__8819\ : CascadeMux
    port map (
            O => \N__42772\,
            I => \N__42737\
        );

    \I__8818\ : CascadeMux
    port map (
            O => \N__42771\,
            I => \N__42734\
        );

    \I__8817\ : CascadeMux
    port map (
            O => \N__42770\,
            I => \N__42731\
        );

    \I__8816\ : CascadeMux
    port map (
            O => \N__42769\,
            I => \N__42728\
        );

    \I__8815\ : CascadeMux
    port map (
            O => \N__42768\,
            I => \N__42725\
        );

    \I__8814\ : CascadeMux
    port map (
            O => \N__42767\,
            I => \N__42722\
        );

    \I__8813\ : CascadeMux
    port map (
            O => \N__42766\,
            I => \N__42719\
        );

    \I__8812\ : CascadeMux
    port map (
            O => \N__42765\,
            I => \N__42716\
        );

    \I__8811\ : CascadeMux
    port map (
            O => \N__42764\,
            I => \N__42713\
        );

    \I__8810\ : InMux
    port map (
            O => \N__42763\,
            I => \N__42698\
        );

    \I__8809\ : InMux
    port map (
            O => \N__42762\,
            I => \N__42698\
        );

    \I__8808\ : InMux
    port map (
            O => \N__42761\,
            I => \N__42695\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__42758\,
            I => \N__42692\
        );

    \I__8806\ : InMux
    port map (
            O => \N__42755\,
            I => \N__42685\
        );

    \I__8805\ : InMux
    port map (
            O => \N__42752\,
            I => \N__42685\
        );

    \I__8804\ : InMux
    port map (
            O => \N__42749\,
            I => \N__42685\
        );

    \I__8803\ : InMux
    port map (
            O => \N__42746\,
            I => \N__42676\
        );

    \I__8802\ : InMux
    port map (
            O => \N__42743\,
            I => \N__42676\
        );

    \I__8801\ : InMux
    port map (
            O => \N__42740\,
            I => \N__42676\
        );

    \I__8800\ : InMux
    port map (
            O => \N__42737\,
            I => \N__42676\
        );

    \I__8799\ : InMux
    port map (
            O => \N__42734\,
            I => \N__42667\
        );

    \I__8798\ : InMux
    port map (
            O => \N__42731\,
            I => \N__42667\
        );

    \I__8797\ : InMux
    port map (
            O => \N__42728\,
            I => \N__42667\
        );

    \I__8796\ : InMux
    port map (
            O => \N__42725\,
            I => \N__42667\
        );

    \I__8795\ : InMux
    port map (
            O => \N__42722\,
            I => \N__42658\
        );

    \I__8794\ : InMux
    port map (
            O => \N__42719\,
            I => \N__42658\
        );

    \I__8793\ : InMux
    port map (
            O => \N__42716\,
            I => \N__42658\
        );

    \I__8792\ : InMux
    port map (
            O => \N__42713\,
            I => \N__42658\
        );

    \I__8791\ : CascadeMux
    port map (
            O => \N__42712\,
            I => \N__42655\
        );

    \I__8790\ : CascadeMux
    port map (
            O => \N__42711\,
            I => \N__42652\
        );

    \I__8789\ : CascadeMux
    port map (
            O => \N__42710\,
            I => \N__42649\
        );

    \I__8788\ : CascadeMux
    port map (
            O => \N__42709\,
            I => \N__42646\
        );

    \I__8787\ : CascadeMux
    port map (
            O => \N__42708\,
            I => \N__42643\
        );

    \I__8786\ : CascadeMux
    port map (
            O => \N__42707\,
            I => \N__42640\
        );

    \I__8785\ : CascadeMux
    port map (
            O => \N__42706\,
            I => \N__42637\
        );

    \I__8784\ : CascadeMux
    port map (
            O => \N__42705\,
            I => \N__42634\
        );

    \I__8783\ : InMux
    port map (
            O => \N__42704\,
            I => \N__42627\
        );

    \I__8782\ : CascadeMux
    port map (
            O => \N__42703\,
            I => \N__42624\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__42698\,
            I => \N__42608\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__42695\,
            I => \N__42608\
        );

    \I__8779\ : Span4Mux_s1_h
    port map (
            O => \N__42692\,
            I => \N__42602\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__42685\,
            I => \N__42586\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__42676\,
            I => \N__42586\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__42667\,
            I => \N__42586\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__42658\,
            I => \N__42586\
        );

    \I__8774\ : InMux
    port map (
            O => \N__42655\,
            I => \N__42577\
        );

    \I__8773\ : InMux
    port map (
            O => \N__42652\,
            I => \N__42577\
        );

    \I__8772\ : InMux
    port map (
            O => \N__42649\,
            I => \N__42577\
        );

    \I__8771\ : InMux
    port map (
            O => \N__42646\,
            I => \N__42577\
        );

    \I__8770\ : InMux
    port map (
            O => \N__42643\,
            I => \N__42568\
        );

    \I__8769\ : InMux
    port map (
            O => \N__42640\,
            I => \N__42568\
        );

    \I__8768\ : InMux
    port map (
            O => \N__42637\,
            I => \N__42568\
        );

    \I__8767\ : InMux
    port map (
            O => \N__42634\,
            I => \N__42568\
        );

    \I__8766\ : CascadeMux
    port map (
            O => \N__42633\,
            I => \N__42565\
        );

    \I__8765\ : CascadeMux
    port map (
            O => \N__42632\,
            I => \N__42562\
        );

    \I__8764\ : CascadeMux
    port map (
            O => \N__42631\,
            I => \N__42559\
        );

    \I__8763\ : CascadeMux
    port map (
            O => \N__42630\,
            I => \N__42556\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__42627\,
            I => \N__42553\
        );

    \I__8761\ : InMux
    port map (
            O => \N__42624\,
            I => \N__42546\
        );

    \I__8760\ : CascadeMux
    port map (
            O => \N__42623\,
            I => \N__42543\
        );

    \I__8759\ : CascadeMux
    port map (
            O => \N__42622\,
            I => \N__42539\
        );

    \I__8758\ : CascadeMux
    port map (
            O => \N__42621\,
            I => \N__42535\
        );

    \I__8757\ : CascadeMux
    port map (
            O => \N__42620\,
            I => \N__42531\
        );

    \I__8756\ : CascadeMux
    port map (
            O => \N__42619\,
            I => \N__42527\
        );

    \I__8755\ : CascadeMux
    port map (
            O => \N__42618\,
            I => \N__42523\
        );

    \I__8754\ : CascadeMux
    port map (
            O => \N__42617\,
            I => \N__42519\
        );

    \I__8753\ : CascadeMux
    port map (
            O => \N__42616\,
            I => \N__42515\
        );

    \I__8752\ : CascadeMux
    port map (
            O => \N__42615\,
            I => \N__42510\
        );

    \I__8751\ : CascadeMux
    port map (
            O => \N__42614\,
            I => \N__42506\
        );

    \I__8750\ : CascadeMux
    port map (
            O => \N__42613\,
            I => \N__42502\
        );

    \I__8749\ : Span4Mux_s2_h
    port map (
            O => \N__42608\,
            I => \N__42498\
        );

    \I__8748\ : InMux
    port map (
            O => \N__42607\,
            I => \N__42493\
        );

    \I__8747\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42493\
        );

    \I__8746\ : InMux
    port map (
            O => \N__42605\,
            I => \N__42490\
        );

    \I__8745\ : Span4Mux_h
    port map (
            O => \N__42602\,
            I => \N__42477\
        );

    \I__8744\ : CascadeMux
    port map (
            O => \N__42601\,
            I => \N__42474\
        );

    \I__8743\ : CascadeMux
    port map (
            O => \N__42600\,
            I => \N__42471\
        );

    \I__8742\ : CascadeMux
    port map (
            O => \N__42599\,
            I => \N__42468\
        );

    \I__8741\ : CascadeMux
    port map (
            O => \N__42598\,
            I => \N__42465\
        );

    \I__8740\ : CascadeMux
    port map (
            O => \N__42597\,
            I => \N__42462\
        );

    \I__8739\ : CascadeMux
    port map (
            O => \N__42596\,
            I => \N__42459\
        );

    \I__8738\ : CascadeMux
    port map (
            O => \N__42595\,
            I => \N__42456\
        );

    \I__8737\ : Span4Mux_v
    port map (
            O => \N__42586\,
            I => \N__42445\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__42577\,
            I => \N__42445\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__42568\,
            I => \N__42445\
        );

    \I__8734\ : InMux
    port map (
            O => \N__42565\,
            I => \N__42440\
        );

    \I__8733\ : InMux
    port map (
            O => \N__42562\,
            I => \N__42440\
        );

    \I__8732\ : InMux
    port map (
            O => \N__42559\,
            I => \N__42435\
        );

    \I__8731\ : InMux
    port map (
            O => \N__42556\,
            I => \N__42435\
        );

    \I__8730\ : Span4Mux_s1_h
    port map (
            O => \N__42553\,
            I => \N__42432\
        );

    \I__8729\ : InMux
    port map (
            O => \N__42552\,
            I => \N__42429\
        );

    \I__8728\ : CascadeMux
    port map (
            O => \N__42551\,
            I => \N__42425\
        );

    \I__8727\ : CascadeMux
    port map (
            O => \N__42550\,
            I => \N__42421\
        );

    \I__8726\ : CascadeMux
    port map (
            O => \N__42549\,
            I => \N__42417\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__42546\,
            I => \N__42413\
        );

    \I__8724\ : InMux
    port map (
            O => \N__42543\,
            I => \N__42396\
        );

    \I__8723\ : InMux
    port map (
            O => \N__42542\,
            I => \N__42396\
        );

    \I__8722\ : InMux
    port map (
            O => \N__42539\,
            I => \N__42396\
        );

    \I__8721\ : InMux
    port map (
            O => \N__42538\,
            I => \N__42396\
        );

    \I__8720\ : InMux
    port map (
            O => \N__42535\,
            I => \N__42396\
        );

    \I__8719\ : InMux
    port map (
            O => \N__42534\,
            I => \N__42396\
        );

    \I__8718\ : InMux
    port map (
            O => \N__42531\,
            I => \N__42396\
        );

    \I__8717\ : InMux
    port map (
            O => \N__42530\,
            I => \N__42396\
        );

    \I__8716\ : InMux
    port map (
            O => \N__42527\,
            I => \N__42379\
        );

    \I__8715\ : InMux
    port map (
            O => \N__42526\,
            I => \N__42379\
        );

    \I__8714\ : InMux
    port map (
            O => \N__42523\,
            I => \N__42379\
        );

    \I__8713\ : InMux
    port map (
            O => \N__42522\,
            I => \N__42379\
        );

    \I__8712\ : InMux
    port map (
            O => \N__42519\,
            I => \N__42379\
        );

    \I__8711\ : InMux
    port map (
            O => \N__42518\,
            I => \N__42379\
        );

    \I__8710\ : InMux
    port map (
            O => \N__42515\,
            I => \N__42379\
        );

    \I__8709\ : InMux
    port map (
            O => \N__42514\,
            I => \N__42379\
        );

    \I__8708\ : InMux
    port map (
            O => \N__42513\,
            I => \N__42364\
        );

    \I__8707\ : InMux
    port map (
            O => \N__42510\,
            I => \N__42364\
        );

    \I__8706\ : InMux
    port map (
            O => \N__42509\,
            I => \N__42364\
        );

    \I__8705\ : InMux
    port map (
            O => \N__42506\,
            I => \N__42364\
        );

    \I__8704\ : InMux
    port map (
            O => \N__42505\,
            I => \N__42364\
        );

    \I__8703\ : InMux
    port map (
            O => \N__42502\,
            I => \N__42364\
        );

    \I__8702\ : InMux
    port map (
            O => \N__42501\,
            I => \N__42364\
        );

    \I__8701\ : Span4Mux_v
    port map (
            O => \N__42498\,
            I => \N__42353\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__42493\,
            I => \N__42348\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__42490\,
            I => \N__42348\
        );

    \I__8698\ : InMux
    port map (
            O => \N__42489\,
            I => \N__42339\
        );

    \I__8697\ : InMux
    port map (
            O => \N__42488\,
            I => \N__42330\
        );

    \I__8696\ : InMux
    port map (
            O => \N__42487\,
            I => \N__42330\
        );

    \I__8695\ : InMux
    port map (
            O => \N__42486\,
            I => \N__42330\
        );

    \I__8694\ : InMux
    port map (
            O => \N__42485\,
            I => \N__42330\
        );

    \I__8693\ : InMux
    port map (
            O => \N__42484\,
            I => \N__42319\
        );

    \I__8692\ : InMux
    port map (
            O => \N__42483\,
            I => \N__42319\
        );

    \I__8691\ : InMux
    port map (
            O => \N__42482\,
            I => \N__42319\
        );

    \I__8690\ : InMux
    port map (
            O => \N__42481\,
            I => \N__42319\
        );

    \I__8689\ : InMux
    port map (
            O => \N__42480\,
            I => \N__42319\
        );

    \I__8688\ : Span4Mux_h
    port map (
            O => \N__42477\,
            I => \N__42316\
        );

    \I__8687\ : InMux
    port map (
            O => \N__42474\,
            I => \N__42309\
        );

    \I__8686\ : InMux
    port map (
            O => \N__42471\,
            I => \N__42309\
        );

    \I__8685\ : InMux
    port map (
            O => \N__42468\,
            I => \N__42309\
        );

    \I__8684\ : InMux
    port map (
            O => \N__42465\,
            I => \N__42300\
        );

    \I__8683\ : InMux
    port map (
            O => \N__42462\,
            I => \N__42300\
        );

    \I__8682\ : InMux
    port map (
            O => \N__42459\,
            I => \N__42300\
        );

    \I__8681\ : InMux
    port map (
            O => \N__42456\,
            I => \N__42300\
        );

    \I__8680\ : CascadeMux
    port map (
            O => \N__42455\,
            I => \N__42297\
        );

    \I__8679\ : CascadeMux
    port map (
            O => \N__42454\,
            I => \N__42294\
        );

    \I__8678\ : CascadeMux
    port map (
            O => \N__42453\,
            I => \N__42291\
        );

    \I__8677\ : CascadeMux
    port map (
            O => \N__42452\,
            I => \N__42288\
        );

    \I__8676\ : Span4Mux_h
    port map (
            O => \N__42445\,
            I => \N__42281\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__42440\,
            I => \N__42281\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__42435\,
            I => \N__42281\
        );

    \I__8673\ : Span4Mux_h
    port map (
            O => \N__42432\,
            I => \N__42278\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__42429\,
            I => \N__42275\
        );

    \I__8671\ : InMux
    port map (
            O => \N__42428\,
            I => \N__42260\
        );

    \I__8670\ : InMux
    port map (
            O => \N__42425\,
            I => \N__42260\
        );

    \I__8669\ : InMux
    port map (
            O => \N__42424\,
            I => \N__42260\
        );

    \I__8668\ : InMux
    port map (
            O => \N__42421\,
            I => \N__42260\
        );

    \I__8667\ : InMux
    port map (
            O => \N__42420\,
            I => \N__42260\
        );

    \I__8666\ : InMux
    port map (
            O => \N__42417\,
            I => \N__42260\
        );

    \I__8665\ : InMux
    port map (
            O => \N__42416\,
            I => \N__42260\
        );

    \I__8664\ : Span4Mux_v
    port map (
            O => \N__42413\,
            I => \N__42251\
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__42396\,
            I => \N__42251\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__42379\,
            I => \N__42251\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__42364\,
            I => \N__42251\
        );

    \I__8660\ : CascadeMux
    port map (
            O => \N__42363\,
            I => \N__42248\
        );

    \I__8659\ : CascadeMux
    port map (
            O => \N__42362\,
            I => \N__42245\
        );

    \I__8658\ : CascadeMux
    port map (
            O => \N__42361\,
            I => \N__42242\
        );

    \I__8657\ : CascadeMux
    port map (
            O => \N__42360\,
            I => \N__42239\
        );

    \I__8656\ : CascadeMux
    port map (
            O => \N__42359\,
            I => \N__42236\
        );

    \I__8655\ : CascadeMux
    port map (
            O => \N__42358\,
            I => \N__42233\
        );

    \I__8654\ : CascadeMux
    port map (
            O => \N__42357\,
            I => \N__42230\
        );

    \I__8653\ : CascadeMux
    port map (
            O => \N__42356\,
            I => \N__42227\
        );

    \I__8652\ : Span4Mux_v
    port map (
            O => \N__42353\,
            I => \N__42213\
        );

    \I__8651\ : Span4Mux_s2_h
    port map (
            O => \N__42348\,
            I => \N__42213\
        );

    \I__8650\ : InMux
    port map (
            O => \N__42347\,
            I => \N__42206\
        );

    \I__8649\ : InMux
    port map (
            O => \N__42346\,
            I => \N__42206\
        );

    \I__8648\ : InMux
    port map (
            O => \N__42345\,
            I => \N__42203\
        );

    \I__8647\ : CascadeMux
    port map (
            O => \N__42344\,
            I => \N__42199\
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__42343\,
            I => \N__42195\
        );

    \I__8645\ : CascadeMux
    port map (
            O => \N__42342\,
            I => \N__42191\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__42339\,
            I => \N__42182\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__42330\,
            I => \N__42182\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__42319\,
            I => \N__42182\
        );

    \I__8641\ : Span4Mux_h
    port map (
            O => \N__42316\,
            I => \N__42179\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__42309\,
            I => \N__42174\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__42300\,
            I => \N__42174\
        );

    \I__8638\ : InMux
    port map (
            O => \N__42297\,
            I => \N__42165\
        );

    \I__8637\ : InMux
    port map (
            O => \N__42294\,
            I => \N__42165\
        );

    \I__8636\ : InMux
    port map (
            O => \N__42291\,
            I => \N__42165\
        );

    \I__8635\ : InMux
    port map (
            O => \N__42288\,
            I => \N__42165\
        );

    \I__8634\ : Span4Mux_v
    port map (
            O => \N__42281\,
            I => \N__42162\
        );

    \I__8633\ : Span4Mux_h
    port map (
            O => \N__42278\,
            I => \N__42153\
        );

    \I__8632\ : Span4Mux_v
    port map (
            O => \N__42275\,
            I => \N__42153\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__42260\,
            I => \N__42153\
        );

    \I__8630\ : Span4Mux_v
    port map (
            O => \N__42251\,
            I => \N__42153\
        );

    \I__8629\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42144\
        );

    \I__8628\ : InMux
    port map (
            O => \N__42245\,
            I => \N__42144\
        );

    \I__8627\ : InMux
    port map (
            O => \N__42242\,
            I => \N__42144\
        );

    \I__8626\ : InMux
    port map (
            O => \N__42239\,
            I => \N__42144\
        );

    \I__8625\ : InMux
    port map (
            O => \N__42236\,
            I => \N__42135\
        );

    \I__8624\ : InMux
    port map (
            O => \N__42233\,
            I => \N__42135\
        );

    \I__8623\ : InMux
    port map (
            O => \N__42230\,
            I => \N__42135\
        );

    \I__8622\ : InMux
    port map (
            O => \N__42227\,
            I => \N__42135\
        );

    \I__8621\ : CascadeMux
    port map (
            O => \N__42226\,
            I => \N__42132\
        );

    \I__8620\ : CascadeMux
    port map (
            O => \N__42225\,
            I => \N__42129\
        );

    \I__8619\ : CascadeMux
    port map (
            O => \N__42224\,
            I => \N__42126\
        );

    \I__8618\ : CascadeMux
    port map (
            O => \N__42223\,
            I => \N__42123\
        );

    \I__8617\ : CascadeMux
    port map (
            O => \N__42222\,
            I => \N__42120\
        );

    \I__8616\ : CascadeMux
    port map (
            O => \N__42221\,
            I => \N__42117\
        );

    \I__8615\ : CascadeMux
    port map (
            O => \N__42220\,
            I => \N__42114\
        );

    \I__8614\ : CascadeMux
    port map (
            O => \N__42219\,
            I => \N__42111\
        );

    \I__8613\ : InMux
    port map (
            O => \N__42218\,
            I => \N__42107\
        );

    \I__8612\ : Span4Mux_h
    port map (
            O => \N__42213\,
            I => \N__42103\
        );

    \I__8611\ : InMux
    port map (
            O => \N__42212\,
            I => \N__42100\
        );

    \I__8610\ : InMux
    port map (
            O => \N__42211\,
            I => \N__42092\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__42206\,
            I => \N__42086\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__42203\,
            I => \N__42086\
        );

    \I__8607\ : InMux
    port map (
            O => \N__42202\,
            I => \N__42071\
        );

    \I__8606\ : InMux
    port map (
            O => \N__42199\,
            I => \N__42071\
        );

    \I__8605\ : InMux
    port map (
            O => \N__42198\,
            I => \N__42071\
        );

    \I__8604\ : InMux
    port map (
            O => \N__42195\,
            I => \N__42071\
        );

    \I__8603\ : InMux
    port map (
            O => \N__42194\,
            I => \N__42071\
        );

    \I__8602\ : InMux
    port map (
            O => \N__42191\,
            I => \N__42071\
        );

    \I__8601\ : InMux
    port map (
            O => \N__42190\,
            I => \N__42071\
        );

    \I__8600\ : CascadeMux
    port map (
            O => \N__42189\,
            I => \N__42068\
        );

    \I__8599\ : Span4Mux_v
    port map (
            O => \N__42182\,
            I => \N__42065\
        );

    \I__8598\ : Span4Mux_h
    port map (
            O => \N__42179\,
            I => \N__42062\
        );

    \I__8597\ : Span4Mux_v
    port map (
            O => \N__42174\,
            I => \N__42057\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__42165\,
            I => \N__42057\
        );

    \I__8595\ : Span4Mux_v
    port map (
            O => \N__42162\,
            I => \N__42048\
        );

    \I__8594\ : Span4Mux_h
    port map (
            O => \N__42153\,
            I => \N__42048\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__42144\,
            I => \N__42048\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__42135\,
            I => \N__42048\
        );

    \I__8591\ : InMux
    port map (
            O => \N__42132\,
            I => \N__42039\
        );

    \I__8590\ : InMux
    port map (
            O => \N__42129\,
            I => \N__42039\
        );

    \I__8589\ : InMux
    port map (
            O => \N__42126\,
            I => \N__42039\
        );

    \I__8588\ : InMux
    port map (
            O => \N__42123\,
            I => \N__42039\
        );

    \I__8587\ : InMux
    port map (
            O => \N__42120\,
            I => \N__42034\
        );

    \I__8586\ : InMux
    port map (
            O => \N__42117\,
            I => \N__42034\
        );

    \I__8585\ : InMux
    port map (
            O => \N__42114\,
            I => \N__42029\
        );

    \I__8584\ : InMux
    port map (
            O => \N__42111\,
            I => \N__42029\
        );

    \I__8583\ : InMux
    port map (
            O => \N__42110\,
            I => \N__42026\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__42107\,
            I => \N__42023\
        );

    \I__8581\ : InMux
    port map (
            O => \N__42106\,
            I => \N__42020\
        );

    \I__8580\ : Span4Mux_h
    port map (
            O => \N__42103\,
            I => \N__42016\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__42100\,
            I => \N__42013\
        );

    \I__8578\ : InMux
    port map (
            O => \N__42099\,
            I => \N__42008\
        );

    \I__8577\ : InMux
    port map (
            O => \N__42098\,
            I => \N__42008\
        );

    \I__8576\ : InMux
    port map (
            O => \N__42097\,
            I => \N__42005\
        );

    \I__8575\ : CascadeMux
    port map (
            O => \N__42096\,
            I => \N__41993\
        );

    \I__8574\ : CascadeMux
    port map (
            O => \N__42095\,
            I => \N__41990\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__42092\,
            I => \N__41986\
        );

    \I__8572\ : InMux
    port map (
            O => \N__42091\,
            I => \N__41983\
        );

    \I__8571\ : Span4Mux_s3_h
    port map (
            O => \N__42086\,
            I => \N__41980\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__42071\,
            I => \N__41977\
        );

    \I__8569\ : InMux
    port map (
            O => \N__42068\,
            I => \N__41974\
        );

    \I__8568\ : Span4Mux_v
    port map (
            O => \N__42065\,
            I => \N__41971\
        );

    \I__8567\ : Span4Mux_v
    port map (
            O => \N__42062\,
            I => \N__41966\
        );

    \I__8566\ : Span4Mux_v
    port map (
            O => \N__42057\,
            I => \N__41966\
        );

    \I__8565\ : Span4Mux_h
    port map (
            O => \N__42048\,
            I => \N__41957\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__42039\,
            I => \N__41957\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__42034\,
            I => \N__41957\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__42029\,
            I => \N__41957\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__42026\,
            I => \N__41950\
        );

    \I__8560\ : Span4Mux_s1_v
    port map (
            O => \N__42023\,
            I => \N__41950\
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__42020\,
            I => \N__41950\
        );

    \I__8558\ : InMux
    port map (
            O => \N__42019\,
            I => \N__41947\
        );

    \I__8557\ : Span4Mux_h
    port map (
            O => \N__42016\,
            I => \N__41944\
        );

    \I__8556\ : Span4Mux_s3_h
    port map (
            O => \N__42013\,
            I => \N__41941\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__42008\,
            I => \N__41936\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__42005\,
            I => \N__41936\
        );

    \I__8553\ : InMux
    port map (
            O => \N__42004\,
            I => \N__41927\
        );

    \I__8552\ : InMux
    port map (
            O => \N__42003\,
            I => \N__41927\
        );

    \I__8551\ : InMux
    port map (
            O => \N__42002\,
            I => \N__41927\
        );

    \I__8550\ : InMux
    port map (
            O => \N__42001\,
            I => \N__41927\
        );

    \I__8549\ : InMux
    port map (
            O => \N__42000\,
            I => \N__41916\
        );

    \I__8548\ : InMux
    port map (
            O => \N__41999\,
            I => \N__41916\
        );

    \I__8547\ : InMux
    port map (
            O => \N__41998\,
            I => \N__41916\
        );

    \I__8546\ : InMux
    port map (
            O => \N__41997\,
            I => \N__41916\
        );

    \I__8545\ : InMux
    port map (
            O => \N__41996\,
            I => \N__41916\
        );

    \I__8544\ : InMux
    port map (
            O => \N__41993\,
            I => \N__41909\
        );

    \I__8543\ : InMux
    port map (
            O => \N__41990\,
            I => \N__41909\
        );

    \I__8542\ : InMux
    port map (
            O => \N__41989\,
            I => \N__41909\
        );

    \I__8541\ : Span12Mux_s10_h
    port map (
            O => \N__41986\,
            I => \N__41906\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__41983\,
            I => \N__41903\
        );

    \I__8539\ : Span4Mux_v
    port map (
            O => \N__41980\,
            I => \N__41896\
        );

    \I__8538\ : Span4Mux_s3_h
    port map (
            O => \N__41977\,
            I => \N__41896\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__41974\,
            I => \N__41896\
        );

    \I__8536\ : Span4Mux_v
    port map (
            O => \N__41971\,
            I => \N__41893\
        );

    \I__8535\ : Span4Mux_v
    port map (
            O => \N__41966\,
            I => \N__41888\
        );

    \I__8534\ : Span4Mux_v
    port map (
            O => \N__41957\,
            I => \N__41888\
        );

    \I__8533\ : Span4Mux_v
    port map (
            O => \N__41950\,
            I => \N__41883\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__41947\,
            I => \N__41883\
        );

    \I__8531\ : Span4Mux_h
    port map (
            O => \N__41944\,
            I => \N__41880\
        );

    \I__8530\ : Span4Mux_v
    port map (
            O => \N__41941\,
            I => \N__41875\
        );

    \I__8529\ : Span4Mux_s3_h
    port map (
            O => \N__41936\,
            I => \N__41875\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__41927\,
            I => \N__41870\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__41916\,
            I => \N__41870\
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__41909\,
            I => \N__41867\
        );

    \I__8525\ : Span12Mux_h
    port map (
            O => \N__41906\,
            I => \N__41864\
        );

    \I__8524\ : Span4Mux_s3_h
    port map (
            O => \N__41903\,
            I => \N__41861\
        );

    \I__8523\ : Span4Mux_v
    port map (
            O => \N__41896\,
            I => \N__41858\
        );

    \I__8522\ : Span4Mux_v
    port map (
            O => \N__41893\,
            I => \N__41851\
        );

    \I__8521\ : Span4Mux_h
    port map (
            O => \N__41888\,
            I => \N__41851\
        );

    \I__8520\ : Span4Mux_v
    port map (
            O => \N__41883\,
            I => \N__41851\
        );

    \I__8519\ : Span4Mux_h
    port map (
            O => \N__41880\,
            I => \N__41842\
        );

    \I__8518\ : Span4Mux_v
    port map (
            O => \N__41875\,
            I => \N__41842\
        );

    \I__8517\ : Span4Mux_s3_h
    port map (
            O => \N__41870\,
            I => \N__41842\
        );

    \I__8516\ : Span4Mux_s3_h
    port map (
            O => \N__41867\,
            I => \N__41842\
        );

    \I__8515\ : Odrv12
    port map (
            O => \N__41864\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8514\ : Odrv4
    port map (
            O => \N__41861\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8513\ : Odrv4
    port map (
            O => \N__41858\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8512\ : Odrv4
    port map (
            O => \N__41851\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8511\ : Odrv4
    port map (
            O => \N__41842\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8510\ : InMux
    port map (
            O => \N__41831\,
            I => \N__41828\
        );

    \I__8509\ : LocalMux
    port map (
            O => \N__41828\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__8508\ : CascadeMux
    port map (
            O => \N__41825\,
            I => \N__41822\
        );

    \I__8507\ : InMux
    port map (
            O => \N__41822\,
            I => \N__41817\
        );

    \I__8506\ : CascadeMux
    port map (
            O => \N__41821\,
            I => \N__41814\
        );

    \I__8505\ : InMux
    port map (
            O => \N__41820\,
            I => \N__41811\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__41817\,
            I => \N__41808\
        );

    \I__8503\ : InMux
    port map (
            O => \N__41814\,
            I => \N__41805\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__41811\,
            I => \N__41802\
        );

    \I__8501\ : Span4Mux_v
    port map (
            O => \N__41808\,
            I => \N__41798\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__41805\,
            I => \N__41795\
        );

    \I__8499\ : Span4Mux_v
    port map (
            O => \N__41802\,
            I => \N__41792\
        );

    \I__8498\ : InMux
    port map (
            O => \N__41801\,
            I => \N__41789\
        );

    \I__8497\ : Odrv4
    port map (
            O => \N__41798\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__8496\ : Odrv12
    port map (
            O => \N__41795\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__8495\ : Odrv4
    port map (
            O => \N__41792\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__41789\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__8493\ : InMux
    port map (
            O => \N__41780\,
            I => \N__41777\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__41777\,
            I => \N__41772\
        );

    \I__8491\ : InMux
    port map (
            O => \N__41776\,
            I => \N__41769\
        );

    \I__8490\ : InMux
    port map (
            O => \N__41775\,
            I => \N__41766\
        );

    \I__8489\ : Span12Mux_s11_h
    port map (
            O => \N__41772\,
            I => \N__41763\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__41769\,
            I => \N__41760\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__41766\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__8486\ : Odrv12
    port map (
            O => \N__41763\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__8485\ : Odrv4
    port map (
            O => \N__41760\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__8484\ : CascadeMux
    port map (
            O => \N__41753\,
            I => \N__41750\
        );

    \I__8483\ : InMux
    port map (
            O => \N__41750\,
            I => \N__41746\
        );

    \I__8482\ : InMux
    port map (
            O => \N__41749\,
            I => \N__41742\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__41746\,
            I => \N__41739\
        );

    \I__8480\ : InMux
    port map (
            O => \N__41745\,
            I => \N__41736\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__41742\,
            I => \N__41733\
        );

    \I__8478\ : Span4Mux_h
    port map (
            O => \N__41739\,
            I => \N__41728\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__41736\,
            I => \N__41728\
        );

    \I__8476\ : Odrv4
    port map (
            O => \N__41733\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__8475\ : Odrv4
    port map (
            O => \N__41728\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__8474\ : CascadeMux
    port map (
            O => \N__41723\,
            I => \N__41719\
        );

    \I__8473\ : CascadeMux
    port map (
            O => \N__41722\,
            I => \N__41715\
        );

    \I__8472\ : InMux
    port map (
            O => \N__41719\,
            I => \N__41712\
        );

    \I__8471\ : InMux
    port map (
            O => \N__41718\,
            I => \N__41709\
        );

    \I__8470\ : InMux
    port map (
            O => \N__41715\,
            I => \N__41706\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__41712\,
            I => \N__41703\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__41709\,
            I => \N__41700\
        );

    \I__8467\ : LocalMux
    port map (
            O => \N__41706\,
            I => \N__41697\
        );

    \I__8466\ : Span4Mux_h
    port map (
            O => \N__41703\,
            I => \N__41691\
        );

    \I__8465\ : Span4Mux_v
    port map (
            O => \N__41700\,
            I => \N__41691\
        );

    \I__8464\ : Span4Mux_v
    port map (
            O => \N__41697\,
            I => \N__41688\
        );

    \I__8463\ : InMux
    port map (
            O => \N__41696\,
            I => \N__41685\
        );

    \I__8462\ : Odrv4
    port map (
            O => \N__41691\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__8461\ : Odrv4
    port map (
            O => \N__41688\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__41685\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__8459\ : CascadeMux
    port map (
            O => \N__41678\,
            I => \N__41675\
        );

    \I__8458\ : InMux
    port map (
            O => \N__41675\,
            I => \N__41671\
        );

    \I__8457\ : InMux
    port map (
            O => \N__41674\,
            I => \N__41667\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__41671\,
            I => \N__41664\
        );

    \I__8455\ : InMux
    port map (
            O => \N__41670\,
            I => \N__41661\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__41667\,
            I => \N__41658\
        );

    \I__8453\ : Span4Mux_v
    port map (
            O => \N__41664\,
            I => \N__41654\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__41661\,
            I => \N__41649\
        );

    \I__8451\ : Sp12to4
    port map (
            O => \N__41658\,
            I => \N__41649\
        );

    \I__8450\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41646\
        );

    \I__8449\ : Odrv4
    port map (
            O => \N__41654\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__8448\ : Odrv12
    port map (
            O => \N__41649\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__41646\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__8446\ : InMux
    port map (
            O => \N__41639\,
            I => \N__41635\
        );

    \I__8445\ : CascadeMux
    port map (
            O => \N__41638\,
            I => \N__41631\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__41635\,
            I => \N__41628\
        );

    \I__8443\ : InMux
    port map (
            O => \N__41634\,
            I => \N__41625\
        );

    \I__8442\ : InMux
    port map (
            O => \N__41631\,
            I => \N__41622\
        );

    \I__8441\ : Span4Mux_h
    port map (
            O => \N__41628\,
            I => \N__41619\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__41625\,
            I => \N__41616\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__41622\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__8438\ : Odrv4
    port map (
            O => \N__41619\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__8437\ : Odrv12
    port map (
            O => \N__41616\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__8436\ : InMux
    port map (
            O => \N__41609\,
            I => \N__41606\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__41606\,
            I => \N__41603\
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__41603\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__8433\ : InMux
    port map (
            O => \N__41600\,
            I => \N__41597\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__41597\,
            I => \N__41594\
        );

    \I__8431\ : Odrv4
    port map (
            O => \N__41594\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__8430\ : CascadeMux
    port map (
            O => \N__41591\,
            I => \N__41588\
        );

    \I__8429\ : InMux
    port map (
            O => \N__41588\,
            I => \N__41585\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__41585\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__8427\ : InMux
    port map (
            O => \N__41582\,
            I => \bfn_16_16_0_\
        );

    \I__8426\ : InMux
    port map (
            O => \N__41579\,
            I => \N__41576\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__41576\,
            I => \N__41573\
        );

    \I__8424\ : Span4Mux_h
    port map (
            O => \N__41573\,
            I => \N__41570\
        );

    \I__8423\ : Odrv4
    port map (
            O => \N__41570\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__8422\ : InMux
    port map (
            O => \N__41567\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__8421\ : CascadeMux
    port map (
            O => \N__41564\,
            I => \N__41561\
        );

    \I__8420\ : InMux
    port map (
            O => \N__41561\,
            I => \N__41558\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__41558\,
            I => \N__41555\
        );

    \I__8418\ : Span4Mux_h
    port map (
            O => \N__41555\,
            I => \N__41552\
        );

    \I__8417\ : Odrv4
    port map (
            O => \N__41552\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__8416\ : InMux
    port map (
            O => \N__41549\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__8415\ : InMux
    port map (
            O => \N__41546\,
            I => \N__41543\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__41543\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__8413\ : InMux
    port map (
            O => \N__41540\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__8412\ : CascadeMux
    port map (
            O => \N__41537\,
            I => \N__41534\
        );

    \I__8411\ : InMux
    port map (
            O => \N__41534\,
            I => \N__41531\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__41531\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__8409\ : InMux
    port map (
            O => \N__41528\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__8408\ : InMux
    port map (
            O => \N__41525\,
            I => \N__41522\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__41522\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__8406\ : InMux
    port map (
            O => \N__41519\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__8405\ : CascadeMux
    port map (
            O => \N__41516\,
            I => \N__41513\
        );

    \I__8404\ : InMux
    port map (
            O => \N__41513\,
            I => \N__41510\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__41510\,
            I => \N__41507\
        );

    \I__8402\ : Span4Mux_h
    port map (
            O => \N__41507\,
            I => \N__41504\
        );

    \I__8401\ : Odrv4
    port map (
            O => \N__41504\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__8400\ : InMux
    port map (
            O => \N__41501\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__8399\ : InMux
    port map (
            O => \N__41498\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__8398\ : InMux
    port map (
            O => \N__41495\,
            I => \N__41492\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__41492\,
            I => \N__41489\
        );

    \I__8396\ : Odrv4
    port map (
            O => \N__41489\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__8395\ : CascadeMux
    port map (
            O => \N__41486\,
            I => \N__41483\
        );

    \I__8394\ : InMux
    port map (
            O => \N__41483\,
            I => \N__41480\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__41480\,
            I => \N__41477\
        );

    \I__8392\ : Span4Mux_h
    port map (
            O => \N__41477\,
            I => \N__41474\
        );

    \I__8391\ : Odrv4
    port map (
            O => \N__41474\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\
        );

    \I__8390\ : InMux
    port map (
            O => \N__41471\,
            I => \bfn_16_15_0_\
        );

    \I__8389\ : InMux
    port map (
            O => \N__41468\,
            I => \N__41465\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__41465\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\
        );

    \I__8387\ : InMux
    port map (
            O => \N__41462\,
            I => \current_shift_inst.un38_control_input_cry_16_s1\
        );

    \I__8386\ : CascadeMux
    port map (
            O => \N__41459\,
            I => \N__41456\
        );

    \I__8385\ : InMux
    port map (
            O => \N__41456\,
            I => \N__41453\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__41453\,
            I => \N__41450\
        );

    \I__8383\ : Odrv4
    port map (
            O => \N__41450\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\
        );

    \I__8382\ : InMux
    port map (
            O => \N__41447\,
            I => \current_shift_inst.un38_control_input_cry_17_s1\
        );

    \I__8381\ : InMux
    port map (
            O => \N__41444\,
            I => \N__41441\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__41441\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\
        );

    \I__8379\ : InMux
    port map (
            O => \N__41438\,
            I => \current_shift_inst.un38_control_input_cry_18_s1\
        );

    \I__8378\ : CascadeMux
    port map (
            O => \N__41435\,
            I => \N__41432\
        );

    \I__8377\ : InMux
    port map (
            O => \N__41432\,
            I => \N__41429\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__41429\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__8375\ : InMux
    port map (
            O => \N__41426\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__8374\ : InMux
    port map (
            O => \N__41423\,
            I => \N__41420\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__41420\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__8372\ : InMux
    port map (
            O => \N__41417\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__8371\ : CascadeMux
    port map (
            O => \N__41414\,
            I => \N__41411\
        );

    \I__8370\ : InMux
    port map (
            O => \N__41411\,
            I => \N__41408\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__41408\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__8368\ : InMux
    port map (
            O => \N__41405\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__8367\ : InMux
    port map (
            O => \N__41402\,
            I => \N__41399\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__41399\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__8365\ : InMux
    port map (
            O => \N__41396\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__8364\ : InMux
    port map (
            O => \N__41393\,
            I => \N__41390\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__41390\,
            I => \N__41387\
        );

    \I__8362\ : Odrv12
    port map (
            O => \N__41387\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\
        );

    \I__8361\ : InMux
    port map (
            O => \N__41384\,
            I => \current_shift_inst.un38_control_input_cry_6_s1\
        );

    \I__8360\ : CascadeMux
    port map (
            O => \N__41381\,
            I => \N__41378\
        );

    \I__8359\ : InMux
    port map (
            O => \N__41378\,
            I => \N__41375\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__41375\,
            I => \N__41372\
        );

    \I__8357\ : Span4Mux_h
    port map (
            O => \N__41372\,
            I => \N__41369\
        );

    \I__8356\ : Span4Mux_v
    port map (
            O => \N__41369\,
            I => \N__41366\
        );

    \I__8355\ : Odrv4
    port map (
            O => \N__41366\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\
        );

    \I__8354\ : InMux
    port map (
            O => \N__41363\,
            I => \bfn_16_14_0_\
        );

    \I__8353\ : InMux
    port map (
            O => \N__41360\,
            I => \N__41357\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__41357\,
            I => \N__41354\
        );

    \I__8351\ : Span4Mux_h
    port map (
            O => \N__41354\,
            I => \N__41351\
        );

    \I__8350\ : Odrv4
    port map (
            O => \N__41351\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\
        );

    \I__8349\ : InMux
    port map (
            O => \N__41348\,
            I => \current_shift_inst.un38_control_input_cry_8_s1\
        );

    \I__8348\ : InMux
    port map (
            O => \N__41345\,
            I => \current_shift_inst.un38_control_input_cry_9_s1\
        );

    \I__8347\ : InMux
    port map (
            O => \N__41342\,
            I => \N__41339\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__41339\,
            I => \N__41336\
        );

    \I__8345\ : Span4Mux_h
    port map (
            O => \N__41336\,
            I => \N__41333\
        );

    \I__8344\ : Odrv4
    port map (
            O => \N__41333\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\
        );

    \I__8343\ : InMux
    port map (
            O => \N__41330\,
            I => \current_shift_inst.un38_control_input_cry_10_s1\
        );

    \I__8342\ : CascadeMux
    port map (
            O => \N__41327\,
            I => \N__41324\
        );

    \I__8341\ : InMux
    port map (
            O => \N__41324\,
            I => \N__41321\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__41321\,
            I => \N__41318\
        );

    \I__8339\ : Span4Mux_h
    port map (
            O => \N__41318\,
            I => \N__41315\
        );

    \I__8338\ : Odrv4
    port map (
            O => \N__41315\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\
        );

    \I__8337\ : InMux
    port map (
            O => \N__41312\,
            I => \current_shift_inst.un38_control_input_cry_11_s1\
        );

    \I__8336\ : InMux
    port map (
            O => \N__41309\,
            I => \N__41306\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__41306\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\
        );

    \I__8334\ : InMux
    port map (
            O => \N__41303\,
            I => \current_shift_inst.un38_control_input_cry_12_s1\
        );

    \I__8333\ : CascadeMux
    port map (
            O => \N__41300\,
            I => \N__41297\
        );

    \I__8332\ : InMux
    port map (
            O => \N__41297\,
            I => \N__41294\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__41294\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\
        );

    \I__8330\ : InMux
    port map (
            O => \N__41291\,
            I => \current_shift_inst.un38_control_input_cry_13_s1\
        );

    \I__8329\ : InMux
    port map (
            O => \N__41288\,
            I => \N__41285\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__41285\,
            I => \N__41282\
        );

    \I__8327\ : Span4Mux_h
    port map (
            O => \N__41282\,
            I => \N__41279\
        );

    \I__8326\ : Odrv4
    port map (
            O => \N__41279\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\
        );

    \I__8325\ : InMux
    port map (
            O => \N__41276\,
            I => \current_shift_inst.un38_control_input_cry_14_s1\
        );

    \I__8324\ : InMux
    port map (
            O => \N__41273\,
            I => \N__41269\
        );

    \I__8323\ : InMux
    port map (
            O => \N__41272\,
            I => \N__41265\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__41269\,
            I => \N__41262\
        );

    \I__8321\ : InMux
    port map (
            O => \N__41268\,
            I => \N__41259\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__41265\,
            I => \N__41256\
        );

    \I__8319\ : Span4Mux_h
    port map (
            O => \N__41262\,
            I => \N__41252\
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__41259\,
            I => \N__41247\
        );

    \I__8317\ : Sp12to4
    port map (
            O => \N__41256\,
            I => \N__41247\
        );

    \I__8316\ : InMux
    port map (
            O => \N__41255\,
            I => \N__41244\
        );

    \I__8315\ : Odrv4
    port map (
            O => \N__41252\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__8314\ : Odrv12
    port map (
            O => \N__41247\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__41244\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__8312\ : InMux
    port map (
            O => \N__41237\,
            I => \N__41234\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__41234\,
            I => \N__41231\
        );

    \I__8310\ : Span4Mux_v
    port map (
            O => \N__41231\,
            I => \N__41228\
        );

    \I__8309\ : Odrv4
    port map (
            O => \N__41228\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__8308\ : CascadeMux
    port map (
            O => \N__41225\,
            I => \N__41222\
        );

    \I__8307\ : InMux
    port map (
            O => \N__41222\,
            I => \N__41219\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__41219\,
            I => \N__41216\
        );

    \I__8305\ : Span4Mux_h
    port map (
            O => \N__41216\,
            I => \N__41213\
        );

    \I__8304\ : Span4Mux_h
    port map (
            O => \N__41213\,
            I => \N__41210\
        );

    \I__8303\ : Odrv4
    port map (
            O => \N__41210\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__8302\ : CascadeMux
    port map (
            O => \N__41207\,
            I => \N__41204\
        );

    \I__8301\ : InMux
    port map (
            O => \N__41204\,
            I => \N__41201\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__41201\,
            I => \N__41198\
        );

    \I__8299\ : Odrv12
    port map (
            O => \N__41198\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__8298\ : InMux
    port map (
            O => \N__41195\,
            I => \current_shift_inst.un38_control_input_cry_2_s1\
        );

    \I__8297\ : CascadeMux
    port map (
            O => \N__41192\,
            I => \N__41189\
        );

    \I__8296\ : InMux
    port map (
            O => \N__41189\,
            I => \N__41186\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__41186\,
            I => \N__41183\
        );

    \I__8294\ : Odrv4
    port map (
            O => \N__41183\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\
        );

    \I__8293\ : InMux
    port map (
            O => \N__41180\,
            I => \current_shift_inst.un38_control_input_cry_3_s1\
        );

    \I__8292\ : InMux
    port map (
            O => \N__41177\,
            I => \N__41174\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__41174\,
            I => \N__41171\
        );

    \I__8290\ : Span4Mux_h
    port map (
            O => \N__41171\,
            I => \N__41168\
        );

    \I__8289\ : Odrv4
    port map (
            O => \N__41168\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\
        );

    \I__8288\ : InMux
    port map (
            O => \N__41165\,
            I => \current_shift_inst.un38_control_input_cry_4_s1\
        );

    \I__8287\ : CascadeMux
    port map (
            O => \N__41162\,
            I => \N__41159\
        );

    \I__8286\ : InMux
    port map (
            O => \N__41159\,
            I => \N__41156\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__41156\,
            I => \N__41153\
        );

    \I__8284\ : Span4Mux_h
    port map (
            O => \N__41153\,
            I => \N__41150\
        );

    \I__8283\ : Span4Mux_h
    port map (
            O => \N__41150\,
            I => \N__41147\
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__41147\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\
        );

    \I__8281\ : InMux
    port map (
            O => \N__41144\,
            I => \current_shift_inst.un38_control_input_cry_5_s1\
        );

    \I__8280\ : InMux
    port map (
            O => \N__41141\,
            I => \N__41137\
        );

    \I__8279\ : InMux
    port map (
            O => \N__41140\,
            I => \N__41134\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__41137\,
            I => \N__41128\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__41134\,
            I => \N__41128\
        );

    \I__8276\ : InMux
    port map (
            O => \N__41133\,
            I => \N__41125\
        );

    \I__8275\ : Span4Mux_h
    port map (
            O => \N__41128\,
            I => \N__41122\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__41125\,
            I => \N__41119\
        );

    \I__8273\ : Span4Mux_v
    port map (
            O => \N__41122\,
            I => \N__41116\
        );

    \I__8272\ : Span12Mux_h
    port map (
            O => \N__41119\,
            I => \N__41113\
        );

    \I__8271\ : Span4Mux_v
    port map (
            O => \N__41116\,
            I => \N__41110\
        );

    \I__8270\ : Odrv12
    port map (
            O => \N__41113\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__8269\ : Odrv4
    port map (
            O => \N__41110\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__8268\ : InMux
    port map (
            O => \N__41105\,
            I => \N__41100\
        );

    \I__8267\ : InMux
    port map (
            O => \N__41104\,
            I => \N__41095\
        );

    \I__8266\ : InMux
    port map (
            O => \N__41103\,
            I => \N__41095\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__41100\,
            I => \N__41089\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__41095\,
            I => \N__41089\
        );

    \I__8263\ : InMux
    port map (
            O => \N__41094\,
            I => \N__41086\
        );

    \I__8262\ : Span12Mux_s11_h
    port map (
            O => \N__41089\,
            I => \N__41083\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__41086\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__8260\ : Odrv12
    port map (
            O => \N__41083\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__8259\ : InMux
    port map (
            O => \N__41078\,
            I => \N__41075\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__41075\,
            I => \N__41069\
        );

    \I__8257\ : InMux
    port map (
            O => \N__41074\,
            I => \N__41066\
        );

    \I__8256\ : InMux
    port map (
            O => \N__41073\,
            I => \N__41063\
        );

    \I__8255\ : InMux
    port map (
            O => \N__41072\,
            I => \N__41060\
        );

    \I__8254\ : Span4Mux_v
    port map (
            O => \N__41069\,
            I => \N__41057\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__41066\,
            I => \N__41054\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__41063\,
            I => \N__41050\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__41060\,
            I => \N__41047\
        );

    \I__8250\ : Sp12to4
    port map (
            O => \N__41057\,
            I => \N__41044\
        );

    \I__8249\ : Span4Mux_v
    port map (
            O => \N__41054\,
            I => \N__41041\
        );

    \I__8248\ : InMux
    port map (
            O => \N__41053\,
            I => \N__41038\
        );

    \I__8247\ : Span4Mux_v
    port map (
            O => \N__41050\,
            I => \N__41035\
        );

    \I__8246\ : Span4Mux_h
    port map (
            O => \N__41047\,
            I => \N__41032\
        );

    \I__8245\ : Odrv12
    port map (
            O => \N__41044\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__8244\ : Odrv4
    port map (
            O => \N__41041\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__41038\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__8242\ : Odrv4
    port map (
            O => \N__41035\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__8241\ : Odrv4
    port map (
            O => \N__41032\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__8240\ : InMux
    port map (
            O => \N__41021\,
            I => \N__41017\
        );

    \I__8239\ : InMux
    port map (
            O => \N__41020\,
            I => \N__41013\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__41017\,
            I => \N__41010\
        );

    \I__8237\ : CascadeMux
    port map (
            O => \N__41016\,
            I => \N__41007\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__41013\,
            I => \N__41004\
        );

    \I__8235\ : Span4Mux_v
    port map (
            O => \N__41010\,
            I => \N__41001\
        );

    \I__8234\ : InMux
    port map (
            O => \N__41007\,
            I => \N__40998\
        );

    \I__8233\ : Span4Mux_v
    port map (
            O => \N__41004\,
            I => \N__40993\
        );

    \I__8232\ : Span4Mux_h
    port map (
            O => \N__41001\,
            I => \N__40993\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__40998\,
            I => \N__40990\
        );

    \I__8230\ : Odrv4
    port map (
            O => \N__40993\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1\
        );

    \I__8229\ : Odrv4
    port map (
            O => \N__40990\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1\
        );

    \I__8228\ : InMux
    port map (
            O => \N__40985\,
            I => \N__40982\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__40982\,
            I => \N__40979\
        );

    \I__8226\ : Span4Mux_h
    port map (
            O => \N__40979\,
            I => \N__40976\
        );

    \I__8225\ : Span4Mux_h
    port map (
            O => \N__40976\,
            I => \N__40973\
        );

    \I__8224\ : Span4Mux_v
    port map (
            O => \N__40973\,
            I => \N__40970\
        );

    \I__8223\ : Odrv4
    port map (
            O => \N__40970\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_0\
        );

    \I__8222\ : CEMux
    port map (
            O => \N__40967\,
            I => \N__40963\
        );

    \I__8221\ : CEMux
    port map (
            O => \N__40966\,
            I => \N__40960\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__40963\,
            I => \N__40957\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__40960\,
            I => \N__40951\
        );

    \I__8218\ : Span4Mux_v
    port map (
            O => \N__40957\,
            I => \N__40948\
        );

    \I__8217\ : CEMux
    port map (
            O => \N__40956\,
            I => \N__40945\
        );

    \I__8216\ : CEMux
    port map (
            O => \N__40955\,
            I => \N__40942\
        );

    \I__8215\ : CEMux
    port map (
            O => \N__40954\,
            I => \N__40938\
        );

    \I__8214\ : Span4Mux_h
    port map (
            O => \N__40951\,
            I => \N__40934\
        );

    \I__8213\ : Span4Mux_v
    port map (
            O => \N__40948\,
            I => \N__40931\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__40945\,
            I => \N__40928\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__40942\,
            I => \N__40925\
        );

    \I__8210\ : CEMux
    port map (
            O => \N__40941\,
            I => \N__40922\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__40938\,
            I => \N__40919\
        );

    \I__8208\ : CEMux
    port map (
            O => \N__40937\,
            I => \N__40916\
        );

    \I__8207\ : Span4Mux_v
    port map (
            O => \N__40934\,
            I => \N__40912\
        );

    \I__8206\ : Span4Mux_h
    port map (
            O => \N__40931\,
            I => \N__40907\
        );

    \I__8205\ : Span4Mux_h
    port map (
            O => \N__40928\,
            I => \N__40907\
        );

    \I__8204\ : Span4Mux_h
    port map (
            O => \N__40925\,
            I => \N__40902\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__40922\,
            I => \N__40902\
        );

    \I__8202\ : Span4Mux_v
    port map (
            O => \N__40919\,
            I => \N__40899\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__40916\,
            I => \N__40896\
        );

    \I__8200\ : CEMux
    port map (
            O => \N__40915\,
            I => \N__40893\
        );

    \I__8199\ : Span4Mux_v
    port map (
            O => \N__40912\,
            I => \N__40888\
        );

    \I__8198\ : Span4Mux_h
    port map (
            O => \N__40907\,
            I => \N__40888\
        );

    \I__8197\ : Span4Mux_h
    port map (
            O => \N__40902\,
            I => \N__40885\
        );

    \I__8196\ : Span4Mux_h
    port map (
            O => \N__40899\,
            I => \N__40878\
        );

    \I__8195\ : Span4Mux_h
    port map (
            O => \N__40896\,
            I => \N__40878\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__40893\,
            I => \N__40878\
        );

    \I__8193\ : Span4Mux_v
    port map (
            O => \N__40888\,
            I => \N__40875\
        );

    \I__8192\ : Span4Mux_v
    port map (
            O => \N__40885\,
            I => \N__40872\
        );

    \I__8191\ : Sp12to4
    port map (
            O => \N__40878\,
            I => \N__40869\
        );

    \I__8190\ : Odrv4
    port map (
            O => \N__40875\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__8189\ : Odrv4
    port map (
            O => \N__40872\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__8188\ : Odrv12
    port map (
            O => \N__40869\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__8187\ : CascadeMux
    port map (
            O => \N__40862\,
            I => \N__40858\
        );

    \I__8186\ : InMux
    port map (
            O => \N__40861\,
            I => \N__40855\
        );

    \I__8185\ : InMux
    port map (
            O => \N__40858\,
            I => \N__40852\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__40855\,
            I => \N__40846\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__40852\,
            I => \N__40846\
        );

    \I__8182\ : InMux
    port map (
            O => \N__40851\,
            I => \N__40842\
        );

    \I__8181\ : Span4Mux_v
    port map (
            O => \N__40846\,
            I => \N__40839\
        );

    \I__8180\ : InMux
    port map (
            O => \N__40845\,
            I => \N__40836\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__40842\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__8178\ : Odrv4
    port map (
            O => \N__40839\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__40836\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__8176\ : InMux
    port map (
            O => \N__40829\,
            I => \N__40826\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__40826\,
            I => \N__40823\
        );

    \I__8174\ : Span4Mux_h
    port map (
            O => \N__40823\,
            I => \N__40820\
        );

    \I__8173\ : Odrv4
    port map (
            O => \N__40820\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__8172\ : InMux
    port map (
            O => \N__40817\,
            I => \N__40814\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__40814\,
            I => \N__40811\
        );

    \I__8170\ : Span4Mux_h
    port map (
            O => \N__40811\,
            I => \N__40808\
        );

    \I__8169\ : Odrv4
    port map (
            O => \N__40808\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__8168\ : InMux
    port map (
            O => \N__40805\,
            I => \N__40801\
        );

    \I__8167\ : CascadeMux
    port map (
            O => \N__40804\,
            I => \N__40798\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__40801\,
            I => \N__40794\
        );

    \I__8165\ : InMux
    port map (
            O => \N__40798\,
            I => \N__40791\
        );

    \I__8164\ : InMux
    port map (
            O => \N__40797\,
            I => \N__40788\
        );

    \I__8163\ : Span4Mux_v
    port map (
            O => \N__40794\,
            I => \N__40783\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__40791\,
            I => \N__40783\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__40788\,
            I => \N__40780\
        );

    \I__8160\ : Span4Mux_v
    port map (
            O => \N__40783\,
            I => \N__40776\
        );

    \I__8159\ : Span4Mux_v
    port map (
            O => \N__40780\,
            I => \N__40773\
        );

    \I__8158\ : InMux
    port map (
            O => \N__40779\,
            I => \N__40770\
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__40776\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__8156\ : Odrv4
    port map (
            O => \N__40773\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__40770\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__8154\ : InMux
    port map (
            O => \N__40763\,
            I => \N__40760\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__40760\,
            I => \N__40757\
        );

    \I__8152\ : Span4Mux_v
    port map (
            O => \N__40757\,
            I => \N__40754\
        );

    \I__8151\ : Odrv4
    port map (
            O => \N__40754\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__8150\ : InMux
    port map (
            O => \N__40751\,
            I => \N__40748\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__40748\,
            I => \N__40745\
        );

    \I__8148\ : Span4Mux_h
    port map (
            O => \N__40745\,
            I => \N__40742\
        );

    \I__8147\ : Odrv4
    port map (
            O => \N__40742\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__8146\ : CascadeMux
    port map (
            O => \N__40739\,
            I => \N__40736\
        );

    \I__8145\ : InMux
    port map (
            O => \N__40736\,
            I => \N__40729\
        );

    \I__8144\ : InMux
    port map (
            O => \N__40735\,
            I => \N__40729\
        );

    \I__8143\ : InMux
    port map (
            O => \N__40734\,
            I => \N__40726\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__40729\,
            I => \N__40721\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__40726\,
            I => \N__40721\
        );

    \I__8140\ : Span4Mux_v
    port map (
            O => \N__40721\,
            I => \N__40717\
        );

    \I__8139\ : InMux
    port map (
            O => \N__40720\,
            I => \N__40714\
        );

    \I__8138\ : Odrv4
    port map (
            O => \N__40717\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__40714\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__8136\ : InMux
    port map (
            O => \N__40709\,
            I => \N__40706\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__40706\,
            I => \N__40703\
        );

    \I__8134\ : Span4Mux_h
    port map (
            O => \N__40703\,
            I => \N__40700\
        );

    \I__8133\ : Odrv4
    port map (
            O => \N__40700\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__8132\ : InMux
    port map (
            O => \N__40697\,
            I => \N__40694\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__40694\,
            I => \N__40691\
        );

    \I__8130\ : Span4Mux_v
    port map (
            O => \N__40691\,
            I => \N__40688\
        );

    \I__8129\ : Odrv4
    port map (
            O => \N__40688\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__8128\ : InMux
    port map (
            O => \N__40685\,
            I => \N__40682\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__40682\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\
        );

    \I__8126\ : InMux
    port map (
            O => \N__40679\,
            I => \N__40676\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__40676\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\
        );

    \I__8124\ : CascadeMux
    port map (
            O => \N__40673\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\
        );

    \I__8123\ : InMux
    port map (
            O => \N__40670\,
            I => \N__40667\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__40667\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\
        );

    \I__8121\ : InMux
    port map (
            O => \N__40664\,
            I => \N__40661\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__40661\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\
        );

    \I__8119\ : CascadeMux
    port map (
            O => \N__40658\,
            I => \N__40655\
        );

    \I__8118\ : InMux
    port map (
            O => \N__40655\,
            I => \N__40652\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__40652\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\
        );

    \I__8116\ : InMux
    port map (
            O => \N__40649\,
            I => \N__40646\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__40646\,
            I => \N__40642\
        );

    \I__8114\ : InMux
    port map (
            O => \N__40645\,
            I => \N__40639\
        );

    \I__8113\ : Span4Mux_h
    port map (
            O => \N__40642\,
            I => \N__40636\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__40639\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__8111\ : Odrv4
    port map (
            O => \N__40636\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__8110\ : InMux
    port map (
            O => \N__40631\,
            I => \N__40611\
        );

    \I__8109\ : InMux
    port map (
            O => \N__40630\,
            I => \N__40611\
        );

    \I__8108\ : InMux
    port map (
            O => \N__40629\,
            I => \N__40599\
        );

    \I__8107\ : InMux
    port map (
            O => \N__40628\,
            I => \N__40599\
        );

    \I__8106\ : InMux
    port map (
            O => \N__40627\,
            I => \N__40594\
        );

    \I__8105\ : InMux
    port map (
            O => \N__40626\,
            I => \N__40594\
        );

    \I__8104\ : InMux
    port map (
            O => \N__40625\,
            I => \N__40589\
        );

    \I__8103\ : InMux
    port map (
            O => \N__40624\,
            I => \N__40589\
        );

    \I__8102\ : InMux
    port map (
            O => \N__40623\,
            I => \N__40584\
        );

    \I__8101\ : InMux
    port map (
            O => \N__40622\,
            I => \N__40584\
        );

    \I__8100\ : InMux
    port map (
            O => \N__40621\,
            I => \N__40568\
        );

    \I__8099\ : InMux
    port map (
            O => \N__40620\,
            I => \N__40568\
        );

    \I__8098\ : InMux
    port map (
            O => \N__40619\,
            I => \N__40568\
        );

    \I__8097\ : InMux
    port map (
            O => \N__40618\,
            I => \N__40568\
        );

    \I__8096\ : InMux
    port map (
            O => \N__40617\,
            I => \N__40563\
        );

    \I__8095\ : InMux
    port map (
            O => \N__40616\,
            I => \N__40563\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__40611\,
            I => \N__40560\
        );

    \I__8093\ : InMux
    port map (
            O => \N__40610\,
            I => \N__40549\
        );

    \I__8092\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40549\
        );

    \I__8091\ : InMux
    port map (
            O => \N__40608\,
            I => \N__40549\
        );

    \I__8090\ : InMux
    port map (
            O => \N__40607\,
            I => \N__40549\
        );

    \I__8089\ : InMux
    port map (
            O => \N__40606\,
            I => \N__40549\
        );

    \I__8088\ : InMux
    port map (
            O => \N__40605\,
            I => \N__40544\
        );

    \I__8087\ : InMux
    port map (
            O => \N__40604\,
            I => \N__40544\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__40599\,
            I => \N__40535\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__40594\,
            I => \N__40535\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__40589\,
            I => \N__40535\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__40584\,
            I => \N__40535\
        );

    \I__8082\ : InMux
    port map (
            O => \N__40583\,
            I => \N__40526\
        );

    \I__8081\ : InMux
    port map (
            O => \N__40582\,
            I => \N__40526\
        );

    \I__8080\ : InMux
    port map (
            O => \N__40581\,
            I => \N__40526\
        );

    \I__8079\ : InMux
    port map (
            O => \N__40580\,
            I => \N__40526\
        );

    \I__8078\ : InMux
    port map (
            O => \N__40579\,
            I => \N__40519\
        );

    \I__8077\ : InMux
    port map (
            O => \N__40578\,
            I => \N__40519\
        );

    \I__8076\ : InMux
    port map (
            O => \N__40577\,
            I => \N__40519\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__40568\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__40563\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8073\ : Odrv4
    port map (
            O => \N__40560\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__40549\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__40544\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8070\ : Odrv4
    port map (
            O => \N__40535\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__40526\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__40519\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8067\ : InMux
    port map (
            O => \N__40502\,
            I => \N__40499\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__40499\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__8065\ : CascadeMux
    port map (
            O => \N__40496\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16_cascade_\
        );

    \I__8064\ : InMux
    port map (
            O => \N__40493\,
            I => \N__40490\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__40490\,
            I => \N__40487\
        );

    \I__8062\ : Span4Mux_h
    port map (
            O => \N__40487\,
            I => \N__40484\
        );

    \I__8061\ : Odrv4
    port map (
            O => \N__40484\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16\
        );

    \I__8060\ : InMux
    port map (
            O => \N__40481\,
            I => \N__40478\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__40478\,
            I => \N__40475\
        );

    \I__8058\ : Sp12to4
    port map (
            O => \N__40475\,
            I => \N__40471\
        );

    \I__8057\ : InMux
    port map (
            O => \N__40474\,
            I => \N__40468\
        );

    \I__8056\ : Span12Mux_s9_h
    port map (
            O => \N__40471\,
            I => \N__40465\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__40468\,
            I => \N__40462\
        );

    \I__8054\ : Span12Mux_v
    port map (
            O => \N__40465\,
            I => \N__40459\
        );

    \I__8053\ : Odrv4
    port map (
            O => \N__40462\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__8052\ : Odrv12
    port map (
            O => \N__40459\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__8051\ : InMux
    port map (
            O => \N__40454\,
            I => \N__40451\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__40451\,
            I => \N__40447\
        );

    \I__8049\ : InMux
    port map (
            O => \N__40450\,
            I => \N__40444\
        );

    \I__8048\ : Span12Mux_s10_h
    port map (
            O => \N__40447\,
            I => \N__40441\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__40444\,
            I => \N__40438\
        );

    \I__8046\ : Span12Mux_v
    port map (
            O => \N__40441\,
            I => \N__40435\
        );

    \I__8045\ : Odrv4
    port map (
            O => \N__40438\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__8044\ : Odrv12
    port map (
            O => \N__40435\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__8043\ : InMux
    port map (
            O => \N__40430\,
            I => \N__40427\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__40427\,
            I => \N__40424\
        );

    \I__8041\ : Odrv4
    port map (
            O => \N__40424\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_31\
        );

    \I__8040\ : InMux
    port map (
            O => \N__40421\,
            I => \N__40418\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__40418\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\
        );

    \I__8038\ : InMux
    port map (
            O => \N__40415\,
            I => \N__40412\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__40412\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\
        );

    \I__8036\ : InMux
    port map (
            O => \N__40409\,
            I => \N__40406\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__40406\,
            I => \N__40403\
        );

    \I__8034\ : Span4Mux_h
    port map (
            O => \N__40403\,
            I => \N__40399\
        );

    \I__8033\ : InMux
    port map (
            O => \N__40402\,
            I => \N__40396\
        );

    \I__8032\ : Odrv4
    port map (
            O => \N__40399\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__40396\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__8030\ : InMux
    port map (
            O => \N__40391\,
            I => \N__40388\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__40388\,
            I => \N__40384\
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__40387\,
            I => \N__40381\
        );

    \I__8027\ : Span4Mux_h
    port map (
            O => \N__40384\,
            I => \N__40378\
        );

    \I__8026\ : InMux
    port map (
            O => \N__40381\,
            I => \N__40375\
        );

    \I__8025\ : Odrv4
    port map (
            O => \N__40378\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__40375\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__8023\ : InMux
    port map (
            O => \N__40370\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_27\
        );

    \I__8022\ : InMux
    port map (
            O => \N__40367\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_28\
        );

    \I__8021\ : InMux
    port map (
            O => \N__40364\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_29\
        );

    \I__8020\ : InMux
    port map (
            O => \N__40361\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_30\
        );

    \I__8019\ : InMux
    port map (
            O => \N__40358\,
            I => \N__40355\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__40355\,
            I => \N__40352\
        );

    \I__8017\ : Span12Mux_s5_h
    port map (
            O => \N__40352\,
            I => \N__40348\
        );

    \I__8016\ : InMux
    port map (
            O => \N__40351\,
            I => \N__40345\
        );

    \I__8015\ : Span12Mux_v
    port map (
            O => \N__40348\,
            I => \N__40342\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__40345\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__8013\ : Odrv12
    port map (
            O => \N__40342\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__8012\ : InMux
    port map (
            O => \N__40337\,
            I => \N__40334\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__40334\,
            I => \N__40331\
        );

    \I__8010\ : Span4Mux_v
    port map (
            O => \N__40331\,
            I => \N__40328\
        );

    \I__8009\ : Sp12to4
    port map (
            O => \N__40328\,
            I => \N__40324\
        );

    \I__8008\ : InMux
    port map (
            O => \N__40327\,
            I => \N__40321\
        );

    \I__8007\ : Span12Mux_s3_h
    port map (
            O => \N__40324\,
            I => \N__40318\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__40321\,
            I => \N__40313\
        );

    \I__8005\ : Span12Mux_h
    port map (
            O => \N__40318\,
            I => \N__40313\
        );

    \I__8004\ : Odrv12
    port map (
            O => \N__40313\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__8003\ : InMux
    port map (
            O => \N__40310\,
            I => \N__40307\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__40307\,
            I => \N__40304\
        );

    \I__8001\ : Span4Mux_s3_h
    port map (
            O => \N__40304\,
            I => \N__40301\
        );

    \I__8000\ : Span4Mux_v
    port map (
            O => \N__40301\,
            I => \N__40297\
        );

    \I__7999\ : InMux
    port map (
            O => \N__40300\,
            I => \N__40294\
        );

    \I__7998\ : Sp12to4
    port map (
            O => \N__40297\,
            I => \N__40291\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__40294\,
            I => \N__40286\
        );

    \I__7996\ : Span12Mux_h
    port map (
            O => \N__40291\,
            I => \N__40286\
        );

    \I__7995\ : Odrv12
    port map (
            O => \N__40286\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__7994\ : InMux
    port map (
            O => \N__40283\,
            I => \N__40280\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__40280\,
            I => \N__40277\
        );

    \I__7992\ : Sp12to4
    port map (
            O => \N__40277\,
            I => \N__40274\
        );

    \I__7991\ : Span12Mux_s6_h
    port map (
            O => \N__40274\,
            I => \N__40270\
        );

    \I__7990\ : InMux
    port map (
            O => \N__40273\,
            I => \N__40267\
        );

    \I__7989\ : Span12Mux_v
    port map (
            O => \N__40270\,
            I => \N__40264\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__40267\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__7987\ : Odrv12
    port map (
            O => \N__40264\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__7986\ : InMux
    port map (
            O => \N__40259\,
            I => \N__40256\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__40256\,
            I => \N__40252\
        );

    \I__7984\ : InMux
    port map (
            O => \N__40255\,
            I => \N__40249\
        );

    \I__7983\ : Span12Mux_s8_h
    port map (
            O => \N__40252\,
            I => \N__40246\
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__40249\,
            I => \N__40243\
        );

    \I__7981\ : Span12Mux_v
    port map (
            O => \N__40246\,
            I => \N__40240\
        );

    \I__7980\ : Odrv4
    port map (
            O => \N__40243\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_27\
        );

    \I__7979\ : Odrv12
    port map (
            O => \N__40240\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_27\
        );

    \I__7978\ : InMux
    port map (
            O => \N__40235\,
            I => \N__40232\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__40232\,
            I => \N__40229\
        );

    \I__7976\ : Span4Mux_h
    port map (
            O => \N__40229\,
            I => \N__40226\
        );

    \I__7975\ : Span4Mux_h
    port map (
            O => \N__40226\,
            I => \N__40222\
        );

    \I__7974\ : InMux
    port map (
            O => \N__40225\,
            I => \N__40219\
        );

    \I__7973\ : Sp12to4
    port map (
            O => \N__40222\,
            I => \N__40216\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__40219\,
            I => \N__40211\
        );

    \I__7971\ : Span12Mux_v
    port map (
            O => \N__40216\,
            I => \N__40211\
        );

    \I__7970\ : Odrv12
    port map (
            O => \N__40211\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__7969\ : InMux
    port map (
            O => \N__40208\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_18\
        );

    \I__7968\ : InMux
    port map (
            O => \N__40205\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_19\
        );

    \I__7967\ : InMux
    port map (
            O => \N__40202\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_20\
        );

    \I__7966\ : InMux
    port map (
            O => \N__40199\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_21\
        );

    \I__7965\ : InMux
    port map (
            O => \N__40196\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_22\
        );

    \I__7964\ : InMux
    port map (
            O => \N__40193\,
            I => \bfn_15_24_0_\
        );

    \I__7963\ : InMux
    port map (
            O => \N__40190\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_24\
        );

    \I__7962\ : InMux
    port map (
            O => \N__40187\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_25\
        );

    \I__7961\ : InMux
    port map (
            O => \N__40184\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_26\
        );

    \I__7960\ : InMux
    port map (
            O => \N__40181\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__7959\ : InMux
    port map (
            O => \N__40178\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__7958\ : InMux
    port map (
            O => \N__40175\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__7957\ : InMux
    port map (
            O => \N__40172\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__7956\ : InMux
    port map (
            O => \N__40169\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__7955\ : InMux
    port map (
            O => \N__40166\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_14\
        );

    \I__7954\ : InMux
    port map (
            O => \N__40163\,
            I => \bfn_15_23_0_\
        );

    \I__7953\ : InMux
    port map (
            O => \N__40160\,
            I => \N__40157\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__40157\,
            I => \N__40153\
        );

    \I__7951\ : InMux
    port map (
            O => \N__40156\,
            I => \N__40150\
        );

    \I__7950\ : Span12Mux_s3_h
    port map (
            O => \N__40153\,
            I => \N__40147\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__40150\,
            I => \N__40144\
        );

    \I__7948\ : Span12Mux_h
    port map (
            O => \N__40147\,
            I => \N__40141\
        );

    \I__7947\ : Odrv4
    port map (
            O => \N__40144\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__7946\ : Odrv12
    port map (
            O => \N__40141\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__7945\ : InMux
    port map (
            O => \N__40136\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_16\
        );

    \I__7944\ : InMux
    port map (
            O => \N__40133\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_17\
        );

    \I__7943\ : InMux
    port map (
            O => \N__40130\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__7942\ : InMux
    port map (
            O => \N__40127\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__7941\ : InMux
    port map (
            O => \N__40124\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__7940\ : InMux
    port map (
            O => \N__40121\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__7939\ : InMux
    port map (
            O => \N__40118\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__7938\ : InMux
    port map (
            O => \N__40115\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__7937\ : InMux
    port map (
            O => \N__40112\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__7936\ : InMux
    port map (
            O => \N__40109\,
            I => \bfn_15_22_0_\
        );

    \I__7935\ : InMux
    port map (
            O => \N__40106\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__7934\ : InMux
    port map (
            O => \N__40103\,
            I => \N__40100\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__40100\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__7932\ : CascadeMux
    port map (
            O => \N__40097\,
            I => \N__40094\
        );

    \I__7931\ : InMux
    port map (
            O => \N__40094\,
            I => \N__40091\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__40091\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__7929\ : InMux
    port map (
            O => \N__40088\,
            I => \N__40085\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__40085\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__7927\ : CascadeMux
    port map (
            O => \N__40082\,
            I => \N__40079\
        );

    \I__7926\ : InMux
    port map (
            O => \N__40079\,
            I => \N__40076\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__40076\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__7924\ : InMux
    port map (
            O => \N__40073\,
            I => \N__40070\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__40070\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__7922\ : CascadeMux
    port map (
            O => \N__40067\,
            I => \N__40064\
        );

    \I__7921\ : InMux
    port map (
            O => \N__40064\,
            I => \N__40061\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__40061\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__7919\ : InMux
    port map (
            O => \N__40058\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__7918\ : InMux
    port map (
            O => \N__40055\,
            I => \N__40052\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__40052\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__7916\ : CascadeMux
    port map (
            O => \N__40049\,
            I => \N__40046\
        );

    \I__7915\ : InMux
    port map (
            O => \N__40046\,
            I => \N__40043\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__40043\,
            I => \N__40040\
        );

    \I__7913\ : Odrv4
    port map (
            O => \N__40040\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__7912\ : InMux
    port map (
            O => \N__40037\,
            I => \N__40034\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__40034\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__7910\ : CascadeMux
    port map (
            O => \N__40031\,
            I => \N__40028\
        );

    \I__7909\ : InMux
    port map (
            O => \N__40028\,
            I => \N__40025\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__40025\,
            I => \N__40022\
        );

    \I__7907\ : Span4Mux_h
    port map (
            O => \N__40022\,
            I => \N__40019\
        );

    \I__7906\ : Span4Mux_v
    port map (
            O => \N__40019\,
            I => \N__40016\
        );

    \I__7905\ : Odrv4
    port map (
            O => \N__40016\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__7904\ : InMux
    port map (
            O => \N__40013\,
            I => \N__40010\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__40010\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__7902\ : CascadeMux
    port map (
            O => \N__40007\,
            I => \N__40004\
        );

    \I__7901\ : InMux
    port map (
            O => \N__40004\,
            I => \N__40001\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__40001\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__7899\ : InMux
    port map (
            O => \N__39998\,
            I => \N__39995\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__39995\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__7897\ : CascadeMux
    port map (
            O => \N__39992\,
            I => \N__39989\
        );

    \I__7896\ : InMux
    port map (
            O => \N__39989\,
            I => \N__39986\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__39986\,
            I => \N__39983\
        );

    \I__7894\ : Span4Mux_v
    port map (
            O => \N__39983\,
            I => \N__39980\
        );

    \I__7893\ : Odrv4
    port map (
            O => \N__39980\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__7892\ : InMux
    port map (
            O => \N__39977\,
            I => \N__39974\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__39974\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__7890\ : CascadeMux
    port map (
            O => \N__39971\,
            I => \N__39968\
        );

    \I__7889\ : InMux
    port map (
            O => \N__39968\,
            I => \N__39965\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__39965\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__7887\ : CascadeMux
    port map (
            O => \N__39962\,
            I => \N__39959\
        );

    \I__7886\ : InMux
    port map (
            O => \N__39959\,
            I => \N__39956\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__39956\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__7884\ : InMux
    port map (
            O => \N__39953\,
            I => \N__39950\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__39950\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__7882\ : CascadeMux
    port map (
            O => \N__39947\,
            I => \N__39944\
        );

    \I__7881\ : InMux
    port map (
            O => \N__39944\,
            I => \N__39941\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__39941\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__7879\ : InMux
    port map (
            O => \N__39938\,
            I => \N__39935\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__39935\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__7877\ : CascadeMux
    port map (
            O => \N__39932\,
            I => \N__39929\
        );

    \I__7876\ : InMux
    port map (
            O => \N__39929\,
            I => \N__39926\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__39926\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__7874\ : InMux
    port map (
            O => \N__39923\,
            I => \N__39920\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__39920\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__7872\ : CascadeMux
    port map (
            O => \N__39917\,
            I => \N__39914\
        );

    \I__7871\ : InMux
    port map (
            O => \N__39914\,
            I => \N__39911\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__39911\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__7869\ : InMux
    port map (
            O => \N__39908\,
            I => \N__39905\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__39905\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__7867\ : InMux
    port map (
            O => \N__39902\,
            I => \N__39898\
        );

    \I__7866\ : InMux
    port map (
            O => \N__39901\,
            I => \N__39894\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__39898\,
            I => \N__39891\
        );

    \I__7864\ : InMux
    port map (
            O => \N__39897\,
            I => \N__39888\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__39894\,
            I => \N__39885\
        );

    \I__7862\ : Span4Mux_v
    port map (
            O => \N__39891\,
            I => \N__39882\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__39888\,
            I => \N__39877\
        );

    \I__7860\ : Span4Mux_v
    port map (
            O => \N__39885\,
            I => \N__39877\
        );

    \I__7859\ : Odrv4
    port map (
            O => \N__39882\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__7858\ : Odrv4
    port map (
            O => \N__39877\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__7857\ : InMux
    port map (
            O => \N__39872\,
            I => \N__39868\
        );

    \I__7856\ : InMux
    port map (
            O => \N__39871\,
            I => \N__39865\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__39868\,
            I => \N__39862\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__39865\,
            I => \N__39859\
        );

    \I__7853\ : Span4Mux_h
    port map (
            O => \N__39862\,
            I => \N__39856\
        );

    \I__7852\ : Span4Mux_h
    port map (
            O => \N__39859\,
            I => \N__39853\
        );

    \I__7851\ : Odrv4
    port map (
            O => \N__39856\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__7850\ : Odrv4
    port map (
            O => \N__39853\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__7849\ : CascadeMux
    port map (
            O => \N__39848\,
            I => \N__39845\
        );

    \I__7848\ : InMux
    port map (
            O => \N__39845\,
            I => \N__39842\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__39842\,
            I => \N__39839\
        );

    \I__7846\ : Odrv4
    port map (
            O => \N__39839\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__7845\ : InMux
    port map (
            O => \N__39836\,
            I => \N__39833\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__39833\,
            I => \N__39830\
        );

    \I__7843\ : Odrv4
    port map (
            O => \N__39830\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__7842\ : CascadeMux
    port map (
            O => \N__39827\,
            I => \N__39824\
        );

    \I__7841\ : InMux
    port map (
            O => \N__39824\,
            I => \N__39821\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__39821\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__7839\ : InMux
    port map (
            O => \N__39818\,
            I => \N__39815\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__39815\,
            I => \N__39812\
        );

    \I__7837\ : Odrv12
    port map (
            O => \N__39812\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__7836\ : CascadeMux
    port map (
            O => \N__39809\,
            I => \N__39806\
        );

    \I__7835\ : InMux
    port map (
            O => \N__39806\,
            I => \N__39803\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__39803\,
            I => \N__39800\
        );

    \I__7833\ : Odrv4
    port map (
            O => \N__39800\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__7832\ : InMux
    port map (
            O => \N__39797\,
            I => \N__39794\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__39794\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__7830\ : CascadeMux
    port map (
            O => \N__39791\,
            I => \N__39788\
        );

    \I__7829\ : InMux
    port map (
            O => \N__39788\,
            I => \N__39785\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__39785\,
            I => \N__39782\
        );

    \I__7827\ : Odrv12
    port map (
            O => \N__39782\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__7826\ : CascadeMux
    port map (
            O => \N__39779\,
            I => \N__39774\
        );

    \I__7825\ : InMux
    port map (
            O => \N__39778\,
            I => \N__39771\
        );

    \I__7824\ : InMux
    port map (
            O => \N__39777\,
            I => \N__39768\
        );

    \I__7823\ : InMux
    port map (
            O => \N__39774\,
            I => \N__39765\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__39771\,
            I => \N__39762\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__39768\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__39765\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__7819\ : Odrv4
    port map (
            O => \N__39762\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__7818\ : InMux
    port map (
            O => \N__39755\,
            I => \N__39750\
        );

    \I__7817\ : InMux
    port map (
            O => \N__39754\,
            I => \N__39747\
        );

    \I__7816\ : InMux
    port map (
            O => \N__39753\,
            I => \N__39744\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__39750\,
            I => \N__39739\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__39747\,
            I => \N__39739\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__39744\,
            I => \N__39733\
        );

    \I__7812\ : Span4Mux_v
    port map (
            O => \N__39739\,
            I => \N__39733\
        );

    \I__7811\ : InMux
    port map (
            O => \N__39738\,
            I => \N__39730\
        );

    \I__7810\ : Odrv4
    port map (
            O => \N__39733\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__39730\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__7808\ : CascadeMux
    port map (
            O => \N__39725\,
            I => \N__39721\
        );

    \I__7807\ : CascadeMux
    port map (
            O => \N__39724\,
            I => \N__39718\
        );

    \I__7806\ : InMux
    port map (
            O => \N__39721\,
            I => \N__39715\
        );

    \I__7805\ : InMux
    port map (
            O => \N__39718\,
            I => \N__39712\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__39715\,
            I => \N__39709\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__39712\,
            I => \N__39703\
        );

    \I__7802\ : Span4Mux_h
    port map (
            O => \N__39709\,
            I => \N__39703\
        );

    \I__7801\ : InMux
    port map (
            O => \N__39708\,
            I => \N__39700\
        );

    \I__7800\ : Span4Mux_v
    port map (
            O => \N__39703\,
            I => \N__39696\
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__39700\,
            I => \N__39693\
        );

    \I__7798\ : InMux
    port map (
            O => \N__39699\,
            I => \N__39690\
        );

    \I__7797\ : Odrv4
    port map (
            O => \N__39696\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__7796\ : Odrv12
    port map (
            O => \N__39693\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__39690\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__7794\ : InMux
    port map (
            O => \N__39683\,
            I => \N__39678\
        );

    \I__7793\ : InMux
    port map (
            O => \N__39682\,
            I => \N__39675\
        );

    \I__7792\ : InMux
    port map (
            O => \N__39681\,
            I => \N__39672\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__39678\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__7790\ : LocalMux
    port map (
            O => \N__39675\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__39672\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__7788\ : CascadeMux
    port map (
            O => \N__39665\,
            I => \N__39661\
        );

    \I__7787\ : InMux
    port map (
            O => \N__39664\,
            I => \N__39643\
        );

    \I__7786\ : InMux
    port map (
            O => \N__39661\,
            I => \N__39643\
        );

    \I__7785\ : InMux
    port map (
            O => \N__39660\,
            I => \N__39640\
        );

    \I__7784\ : InMux
    port map (
            O => \N__39659\,
            I => \N__39628\
        );

    \I__7783\ : InMux
    port map (
            O => \N__39658\,
            I => \N__39628\
        );

    \I__7782\ : InMux
    port map (
            O => \N__39657\,
            I => \N__39615\
        );

    \I__7781\ : InMux
    port map (
            O => \N__39656\,
            I => \N__39615\
        );

    \I__7780\ : InMux
    port map (
            O => \N__39655\,
            I => \N__39615\
        );

    \I__7779\ : InMux
    port map (
            O => \N__39654\,
            I => \N__39615\
        );

    \I__7778\ : InMux
    port map (
            O => \N__39653\,
            I => \N__39615\
        );

    \I__7777\ : InMux
    port map (
            O => \N__39652\,
            I => \N__39615\
        );

    \I__7776\ : InMux
    port map (
            O => \N__39651\,
            I => \N__39606\
        );

    \I__7775\ : InMux
    port map (
            O => \N__39650\,
            I => \N__39606\
        );

    \I__7774\ : InMux
    port map (
            O => \N__39649\,
            I => \N__39606\
        );

    \I__7773\ : InMux
    port map (
            O => \N__39648\,
            I => \N__39606\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__39643\,
            I => \N__39601\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__39640\,
            I => \N__39601\
        );

    \I__7770\ : InMux
    port map (
            O => \N__39639\,
            I => \N__39586\
        );

    \I__7769\ : InMux
    port map (
            O => \N__39638\,
            I => \N__39586\
        );

    \I__7768\ : InMux
    port map (
            O => \N__39637\,
            I => \N__39586\
        );

    \I__7767\ : InMux
    port map (
            O => \N__39636\,
            I => \N__39586\
        );

    \I__7766\ : InMux
    port map (
            O => \N__39635\,
            I => \N__39586\
        );

    \I__7765\ : InMux
    port map (
            O => \N__39634\,
            I => \N__39586\
        );

    \I__7764\ : InMux
    port map (
            O => \N__39633\,
            I => \N__39586\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__39628\,
            I => \N__39582\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__39615\,
            I => \N__39579\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__39606\,
            I => \N__39574\
        );

    \I__7760\ : Span4Mux_v
    port map (
            O => \N__39601\,
            I => \N__39569\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__39586\,
            I => \N__39569\
        );

    \I__7758\ : InMux
    port map (
            O => \N__39585\,
            I => \N__39566\
        );

    \I__7757\ : Span4Mux_v
    port map (
            O => \N__39582\,
            I => \N__39563\
        );

    \I__7756\ : Span4Mux_h
    port map (
            O => \N__39579\,
            I => \N__39560\
        );

    \I__7755\ : InMux
    port map (
            O => \N__39578\,
            I => \N__39555\
        );

    \I__7754\ : InMux
    port map (
            O => \N__39577\,
            I => \N__39555\
        );

    \I__7753\ : Span4Mux_h
    port map (
            O => \N__39574\,
            I => \N__39552\
        );

    \I__7752\ : Odrv4
    port map (
            O => \N__39569\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__39566\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__7750\ : Odrv4
    port map (
            O => \N__39563\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__7749\ : Odrv4
    port map (
            O => \N__39560\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__39555\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__7747\ : Odrv4
    port map (
            O => \N__39552\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__7746\ : CascadeMux
    port map (
            O => \N__39539\,
            I => \N__39534\
        );

    \I__7745\ : InMux
    port map (
            O => \N__39538\,
            I => \N__39531\
        );

    \I__7744\ : InMux
    port map (
            O => \N__39537\,
            I => \N__39528\
        );

    \I__7743\ : InMux
    port map (
            O => \N__39534\,
            I => \N__39525\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__39531\,
            I => \N__39522\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__39528\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__39525\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__7739\ : Odrv4
    port map (
            O => \N__39522\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__7738\ : InMux
    port map (
            O => \N__39515\,
            I => \N__39510\
        );

    \I__7737\ : InMux
    port map (
            O => \N__39514\,
            I => \N__39507\
        );

    \I__7736\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39504\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__39510\,
            I => \N__39501\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__39507\,
            I => \N__39496\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__39504\,
            I => \N__39496\
        );

    \I__7732\ : Span4Mux_v
    port map (
            O => \N__39501\,
            I => \N__39490\
        );

    \I__7731\ : Span4Mux_v
    port map (
            O => \N__39496\,
            I => \N__39490\
        );

    \I__7730\ : InMux
    port map (
            O => \N__39495\,
            I => \N__39487\
        );

    \I__7729\ : Odrv4
    port map (
            O => \N__39490\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__39487\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__7727\ : CascadeMux
    port map (
            O => \N__39482\,
            I => \N__39477\
        );

    \I__7726\ : InMux
    port map (
            O => \N__39481\,
            I => \N__39474\
        );

    \I__7725\ : InMux
    port map (
            O => \N__39480\,
            I => \N__39471\
        );

    \I__7724\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39468\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__39474\,
            I => \N__39463\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__39471\,
            I => \N__39463\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__39468\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__7720\ : Odrv4
    port map (
            O => \N__39463\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__7719\ : InMux
    port map (
            O => \N__39458\,
            I => \N__39455\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__39455\,
            I => \N__39452\
        );

    \I__7717\ : Span4Mux_v
    port map (
            O => \N__39452\,
            I => \N__39447\
        );

    \I__7716\ : InMux
    port map (
            O => \N__39451\,
            I => \N__39444\
        );

    \I__7715\ : InMux
    port map (
            O => \N__39450\,
            I => \N__39441\
        );

    \I__7714\ : Span4Mux_h
    port map (
            O => \N__39447\,
            I => \N__39436\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__39444\,
            I => \N__39436\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__39441\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__7711\ : Odrv4
    port map (
            O => \N__39436\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__7710\ : InMux
    port map (
            O => \N__39431\,
            I => \N__39426\
        );

    \I__7709\ : InMux
    port map (
            O => \N__39430\,
            I => \N__39423\
        );

    \I__7708\ : CascadeMux
    port map (
            O => \N__39429\,
            I => \N__39420\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__39426\,
            I => \N__39414\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__39423\,
            I => \N__39414\
        );

    \I__7705\ : InMux
    port map (
            O => \N__39420\,
            I => \N__39411\
        );

    \I__7704\ : InMux
    port map (
            O => \N__39419\,
            I => \N__39408\
        );

    \I__7703\ : Span4Mux_v
    port map (
            O => \N__39414\,
            I => \N__39405\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__39411\,
            I => \N__39400\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__39408\,
            I => \N__39400\
        );

    \I__7700\ : Span4Mux_v
    port map (
            O => \N__39405\,
            I => \N__39397\
        );

    \I__7699\ : Span4Mux_h
    port map (
            O => \N__39400\,
            I => \N__39394\
        );

    \I__7698\ : Odrv4
    port map (
            O => \N__39397\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__39394\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__7696\ : CascadeMux
    port map (
            O => \N__39389\,
            I => \N__39386\
        );

    \I__7695\ : InMux
    port map (
            O => \N__39386\,
            I => \N__39382\
        );

    \I__7694\ : InMux
    port map (
            O => \N__39385\,
            I => \N__39378\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__39382\,
            I => \N__39375\
        );

    \I__7692\ : InMux
    port map (
            O => \N__39381\,
            I => \N__39372\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__39378\,
            I => \N__39369\
        );

    \I__7690\ : Span4Mux_h
    port map (
            O => \N__39375\,
            I => \N__39364\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__39372\,
            I => \N__39364\
        );

    \I__7688\ : Span4Mux_v
    port map (
            O => \N__39369\,
            I => \N__39358\
        );

    \I__7687\ : Span4Mux_v
    port map (
            O => \N__39364\,
            I => \N__39358\
        );

    \I__7686\ : InMux
    port map (
            O => \N__39363\,
            I => \N__39355\
        );

    \I__7685\ : Odrv4
    port map (
            O => \N__39358\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__39355\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__7683\ : InMux
    port map (
            O => \N__39350\,
            I => \N__39343\
        );

    \I__7682\ : InMux
    port map (
            O => \N__39349\,
            I => \N__39343\
        );

    \I__7681\ : InMux
    port map (
            O => \N__39348\,
            I => \N__39340\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__39343\,
            I => \N__39336\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__39340\,
            I => \N__39333\
        );

    \I__7678\ : InMux
    port map (
            O => \N__39339\,
            I => \N__39330\
        );

    \I__7677\ : Span4Mux_h
    port map (
            O => \N__39336\,
            I => \N__39327\
        );

    \I__7676\ : Sp12to4
    port map (
            O => \N__39333\,
            I => \N__39322\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__39330\,
            I => \N__39322\
        );

    \I__7674\ : Odrv4
    port map (
            O => \N__39327\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__7673\ : Odrv12
    port map (
            O => \N__39322\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__7672\ : InMux
    port map (
            O => \N__39317\,
            I => \N__39314\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__39314\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__7670\ : InMux
    port map (
            O => \N__39311\,
            I => \N__39308\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__39308\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__7668\ : CascadeMux
    port map (
            O => \N__39305\,
            I => \N__39302\
        );

    \I__7667\ : InMux
    port map (
            O => \N__39302\,
            I => \N__39298\
        );

    \I__7666\ : InMux
    port map (
            O => \N__39301\,
            I => \N__39294\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__39298\,
            I => \N__39291\
        );

    \I__7664\ : InMux
    port map (
            O => \N__39297\,
            I => \N__39288\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__39294\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__7662\ : Odrv4
    port map (
            O => \N__39291\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__39288\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__7660\ : InMux
    port map (
            O => \N__39281\,
            I => \N__39276\
        );

    \I__7659\ : InMux
    port map (
            O => \N__39280\,
            I => \N__39273\
        );

    \I__7658\ : InMux
    port map (
            O => \N__39279\,
            I => \N__39270\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__39276\,
            I => \N__39267\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__39273\,
            I => \N__39264\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__39270\,
            I => \N__39260\
        );

    \I__7654\ : Span4Mux_v
    port map (
            O => \N__39267\,
            I => \N__39257\
        );

    \I__7653\ : Span4Mux_v
    port map (
            O => \N__39264\,
            I => \N__39254\
        );

    \I__7652\ : InMux
    port map (
            O => \N__39263\,
            I => \N__39251\
        );

    \I__7651\ : Odrv12
    port map (
            O => \N__39260\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__7650\ : Odrv4
    port map (
            O => \N__39257\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__7649\ : Odrv4
    port map (
            O => \N__39254\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__39251\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__7647\ : CascadeMux
    port map (
            O => \N__39242\,
            I => \N__39237\
        );

    \I__7646\ : InMux
    port map (
            O => \N__39241\,
            I => \N__39234\
        );

    \I__7645\ : InMux
    port map (
            O => \N__39240\,
            I => \N__39231\
        );

    \I__7644\ : InMux
    port map (
            O => \N__39237\,
            I => \N__39228\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__39234\,
            I => \N__39223\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__39231\,
            I => \N__39223\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__39228\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__7640\ : Odrv4
    port map (
            O => \N__39223\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__7639\ : CascadeMux
    port map (
            O => \N__39218\,
            I => \N__39215\
        );

    \I__7638\ : InMux
    port map (
            O => \N__39215\,
            I => \N__39210\
        );

    \I__7637\ : InMux
    port map (
            O => \N__39214\,
            I => \N__39207\
        );

    \I__7636\ : InMux
    port map (
            O => \N__39213\,
            I => \N__39204\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__39210\,
            I => \N__39201\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__39207\,
            I => \N__39198\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__39204\,
            I => \N__39191\
        );

    \I__7632\ : Span4Mux_v
    port map (
            O => \N__39201\,
            I => \N__39191\
        );

    \I__7631\ : Span4Mux_v
    port map (
            O => \N__39198\,
            I => \N__39191\
        );

    \I__7630\ : Span4Mux_v
    port map (
            O => \N__39191\,
            I => \N__39187\
        );

    \I__7629\ : InMux
    port map (
            O => \N__39190\,
            I => \N__39184\
        );

    \I__7628\ : Odrv4
    port map (
            O => \N__39187\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__39184\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__7626\ : InMux
    port map (
            O => \N__39179\,
            I => \N__39175\
        );

    \I__7625\ : CascadeMux
    port map (
            O => \N__39178\,
            I => \N__39171\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__39175\,
            I => \N__39168\
        );

    \I__7623\ : InMux
    port map (
            O => \N__39174\,
            I => \N__39165\
        );

    \I__7622\ : InMux
    port map (
            O => \N__39171\,
            I => \N__39162\
        );

    \I__7621\ : Span4Mux_v
    port map (
            O => \N__39168\,
            I => \N__39159\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__39165\,
            I => \N__39156\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__39162\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__7618\ : Odrv4
    port map (
            O => \N__39159\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__7617\ : Odrv4
    port map (
            O => \N__39156\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__7616\ : InMux
    port map (
            O => \N__39149\,
            I => \N__39144\
        );

    \I__7615\ : InMux
    port map (
            O => \N__39148\,
            I => \N__39141\
        );

    \I__7614\ : InMux
    port map (
            O => \N__39147\,
            I => \N__39138\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__39144\,
            I => \N__39135\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__39141\,
            I => \N__39130\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__39138\,
            I => \N__39130\
        );

    \I__7610\ : Span4Mux_h
    port map (
            O => \N__39135\,
            I => \N__39124\
        );

    \I__7609\ : Span4Mux_v
    port map (
            O => \N__39130\,
            I => \N__39124\
        );

    \I__7608\ : InMux
    port map (
            O => \N__39129\,
            I => \N__39121\
        );

    \I__7607\ : Odrv4
    port map (
            O => \N__39124\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__39121\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__7605\ : InMux
    port map (
            O => \N__39116\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__7604\ : InMux
    port map (
            O => \N__39113\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__7603\ : InMux
    port map (
            O => \N__39110\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__7602\ : InMux
    port map (
            O => \N__39107\,
            I => \N__39104\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__39104\,
            I => \N__39100\
        );

    \I__7600\ : InMux
    port map (
            O => \N__39103\,
            I => \N__39097\
        );

    \I__7599\ : Span4Mux_h
    port map (
            O => \N__39100\,
            I => \N__39093\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__39097\,
            I => \N__39090\
        );

    \I__7597\ : InMux
    port map (
            O => \N__39096\,
            I => \N__39087\
        );

    \I__7596\ : Odrv4
    port map (
            O => \N__39093\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__7595\ : Odrv4
    port map (
            O => \N__39090\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__39087\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__7593\ : CEMux
    port map (
            O => \N__39080\,
            I => \N__39059\
        );

    \I__7592\ : CEMux
    port map (
            O => \N__39079\,
            I => \N__39059\
        );

    \I__7591\ : CEMux
    port map (
            O => \N__39078\,
            I => \N__39059\
        );

    \I__7590\ : CEMux
    port map (
            O => \N__39077\,
            I => \N__39059\
        );

    \I__7589\ : CEMux
    port map (
            O => \N__39076\,
            I => \N__39059\
        );

    \I__7588\ : CEMux
    port map (
            O => \N__39075\,
            I => \N__39059\
        );

    \I__7587\ : CEMux
    port map (
            O => \N__39074\,
            I => \N__39059\
        );

    \I__7586\ : GlobalMux
    port map (
            O => \N__39059\,
            I => \N__39056\
        );

    \I__7585\ : gio2CtrlBuf
    port map (
            O => \N__39056\,
            I => \current_shift_inst.timer_s1.N_163_i_g\
        );

    \I__7584\ : CascadeMux
    port map (
            O => \N__39053\,
            I => \N__39050\
        );

    \I__7583\ : InMux
    port map (
            O => \N__39050\,
            I => \N__39046\
        );

    \I__7582\ : InMux
    port map (
            O => \N__39049\,
            I => \N__39043\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__39046\,
            I => \N__39039\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__39043\,
            I => \N__39036\
        );

    \I__7579\ : InMux
    port map (
            O => \N__39042\,
            I => \N__39033\
        );

    \I__7578\ : Span4Mux_h
    port map (
            O => \N__39039\,
            I => \N__39029\
        );

    \I__7577\ : Span4Mux_h
    port map (
            O => \N__39036\,
            I => \N__39026\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__39033\,
            I => \N__39023\
        );

    \I__7575\ : InMux
    port map (
            O => \N__39032\,
            I => \N__39020\
        );

    \I__7574\ : Odrv4
    port map (
            O => \N__39029\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__7573\ : Odrv4
    port map (
            O => \N__39026\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__7572\ : Odrv12
    port map (
            O => \N__39023\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__39020\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__7570\ : InMux
    port map (
            O => \N__39011\,
            I => \N__39007\
        );

    \I__7569\ : InMux
    port map (
            O => \N__39010\,
            I => \N__39003\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__39007\,
            I => \N__39000\
        );

    \I__7567\ : InMux
    port map (
            O => \N__39006\,
            I => \N__38997\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__39003\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__7565\ : Odrv4
    port map (
            O => \N__39000\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__38997\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__7563\ : InMux
    port map (
            O => \N__38990\,
            I => \N__38983\
        );

    \I__7562\ : InMux
    port map (
            O => \N__38989\,
            I => \N__38983\
        );

    \I__7561\ : InMux
    port map (
            O => \N__38988\,
            I => \N__38980\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__38983\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__38980\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__7558\ : CascadeMux
    port map (
            O => \N__38975\,
            I => \N__38971\
        );

    \I__7557\ : InMux
    port map (
            O => \N__38974\,
            I => \N__38966\
        );

    \I__7556\ : InMux
    port map (
            O => \N__38971\,
            I => \N__38966\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__38966\,
            I => \N__38962\
        );

    \I__7554\ : InMux
    port map (
            O => \N__38965\,
            I => \N__38959\
        );

    \I__7553\ : Span4Mux_v
    port map (
            O => \N__38962\,
            I => \N__38956\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__38959\,
            I => \N__38953\
        );

    \I__7551\ : Span4Mux_h
    port map (
            O => \N__38956\,
            I => \N__38949\
        );

    \I__7550\ : Span4Mux_v
    port map (
            O => \N__38953\,
            I => \N__38946\
        );

    \I__7549\ : InMux
    port map (
            O => \N__38952\,
            I => \N__38943\
        );

    \I__7548\ : Odrv4
    port map (
            O => \N__38949\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__7547\ : Odrv4
    port map (
            O => \N__38946\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__38943\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__7545\ : InMux
    port map (
            O => \N__38936\,
            I => \N__38930\
        );

    \I__7544\ : InMux
    port map (
            O => \N__38935\,
            I => \N__38930\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__38930\,
            I => \N__38926\
        );

    \I__7542\ : InMux
    port map (
            O => \N__38929\,
            I => \N__38923\
        );

    \I__7541\ : Span4Mux_v
    port map (
            O => \N__38926\,
            I => \N__38919\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__38923\,
            I => \N__38916\
        );

    \I__7539\ : InMux
    port map (
            O => \N__38922\,
            I => \N__38913\
        );

    \I__7538\ : Odrv4
    port map (
            O => \N__38919\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__7537\ : Odrv12
    port map (
            O => \N__38916\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__38913\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__7535\ : CascadeMux
    port map (
            O => \N__38906\,
            I => \N__38903\
        );

    \I__7534\ : InMux
    port map (
            O => \N__38903\,
            I => \N__38896\
        );

    \I__7533\ : InMux
    port map (
            O => \N__38902\,
            I => \N__38896\
        );

    \I__7532\ : InMux
    port map (
            O => \N__38901\,
            I => \N__38893\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__38896\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__38893\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__7529\ : InMux
    port map (
            O => \N__38888\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__7528\ : InMux
    port map (
            O => \N__38885\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__7527\ : InMux
    port map (
            O => \N__38882\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__7526\ : InMux
    port map (
            O => \N__38879\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__7525\ : InMux
    port map (
            O => \N__38876\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__7524\ : InMux
    port map (
            O => \N__38873\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__7523\ : InMux
    port map (
            O => \N__38870\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__7522\ : InMux
    port map (
            O => \N__38867\,
            I => \N__38860\
        );

    \I__7521\ : InMux
    port map (
            O => \N__38866\,
            I => \N__38860\
        );

    \I__7520\ : InMux
    port map (
            O => \N__38865\,
            I => \N__38856\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__38860\,
            I => \N__38853\
        );

    \I__7518\ : InMux
    port map (
            O => \N__38859\,
            I => \N__38850\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__38856\,
            I => \N__38847\
        );

    \I__7516\ : Span4Mux_v
    port map (
            O => \N__38853\,
            I => \N__38842\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__38850\,
            I => \N__38842\
        );

    \I__7514\ : Sp12to4
    port map (
            O => \N__38847\,
            I => \N__38839\
        );

    \I__7513\ : Span4Mux_v
    port map (
            O => \N__38842\,
            I => \N__38836\
        );

    \I__7512\ : Odrv12
    port map (
            O => \N__38839\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__7511\ : Odrv4
    port map (
            O => \N__38836\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__7510\ : InMux
    port map (
            O => \N__38831\,
            I => \bfn_15_13_0_\
        );

    \I__7509\ : InMux
    port map (
            O => \N__38828\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__7508\ : InMux
    port map (
            O => \N__38825\,
            I => \bfn_15_11_0_\
        );

    \I__7507\ : CascadeMux
    port map (
            O => \N__38822\,
            I => \N__38818\
        );

    \I__7506\ : CascadeMux
    port map (
            O => \N__38821\,
            I => \N__38815\
        );

    \I__7505\ : InMux
    port map (
            O => \N__38818\,
            I => \N__38812\
        );

    \I__7504\ : InMux
    port map (
            O => \N__38815\,
            I => \N__38809\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__38812\,
            I => \N__38805\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__38809\,
            I => \N__38802\
        );

    \I__7501\ : InMux
    port map (
            O => \N__38808\,
            I => \N__38799\
        );

    \I__7500\ : Span4Mux_h
    port map (
            O => \N__38805\,
            I => \N__38794\
        );

    \I__7499\ : Span4Mux_h
    port map (
            O => \N__38802\,
            I => \N__38794\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__38799\,
            I => \N__38791\
        );

    \I__7497\ : Span4Mux_v
    port map (
            O => \N__38794\,
            I => \N__38787\
        );

    \I__7496\ : Span4Mux_v
    port map (
            O => \N__38791\,
            I => \N__38784\
        );

    \I__7495\ : InMux
    port map (
            O => \N__38790\,
            I => \N__38781\
        );

    \I__7494\ : Odrv4
    port map (
            O => \N__38787\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__7493\ : Odrv4
    port map (
            O => \N__38784\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__38781\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__7491\ : InMux
    port map (
            O => \N__38774\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__7490\ : InMux
    port map (
            O => \N__38771\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__7489\ : InMux
    port map (
            O => \N__38768\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__7488\ : InMux
    port map (
            O => \N__38765\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__7487\ : InMux
    port map (
            O => \N__38762\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__7486\ : CascadeMux
    port map (
            O => \N__38759\,
            I => \N__38756\
        );

    \I__7485\ : InMux
    port map (
            O => \N__38756\,
            I => \N__38753\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__38753\,
            I => \N__38748\
        );

    \I__7483\ : InMux
    port map (
            O => \N__38752\,
            I => \N__38745\
        );

    \I__7482\ : InMux
    port map (
            O => \N__38751\,
            I => \N__38742\
        );

    \I__7481\ : Span4Mux_h
    port map (
            O => \N__38748\,
            I => \N__38737\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__38745\,
            I => \N__38737\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__38742\,
            I => \N__38734\
        );

    \I__7478\ : Span4Mux_v
    port map (
            O => \N__38737\,
            I => \N__38731\
        );

    \I__7477\ : Span4Mux_h
    port map (
            O => \N__38734\,
            I => \N__38727\
        );

    \I__7476\ : Span4Mux_v
    port map (
            O => \N__38731\,
            I => \N__38724\
        );

    \I__7475\ : InMux
    port map (
            O => \N__38730\,
            I => \N__38721\
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__38727\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__7473\ : Odrv4
    port map (
            O => \N__38724\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__38721\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__7471\ : InMux
    port map (
            O => \N__38714\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__7470\ : InMux
    port map (
            O => \N__38711\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__7469\ : InMux
    port map (
            O => \N__38708\,
            I => \bfn_15_12_0_\
        );

    \I__7468\ : InMux
    port map (
            O => \N__38705\,
            I => \N__38701\
        );

    \I__7467\ : InMux
    port map (
            O => \N__38704\,
            I => \N__38698\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__38701\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__38698\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__7464\ : InMux
    port map (
            O => \N__38693\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__7463\ : InMux
    port map (
            O => \N__38690\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__7462\ : InMux
    port map (
            O => \N__38687\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__7461\ : CascadeMux
    port map (
            O => \N__38684\,
            I => \N__38680\
        );

    \I__7460\ : InMux
    port map (
            O => \N__38683\,
            I => \N__38677\
        );

    \I__7459\ : InMux
    port map (
            O => \N__38680\,
            I => \N__38674\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__38677\,
            I => \N__38670\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__38674\,
            I => \N__38667\
        );

    \I__7456\ : InMux
    port map (
            O => \N__38673\,
            I => \N__38664\
        );

    \I__7455\ : Span4Mux_h
    port map (
            O => \N__38670\,
            I => \N__38659\
        );

    \I__7454\ : Span4Mux_h
    port map (
            O => \N__38667\,
            I => \N__38659\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__38664\,
            I => \N__38656\
        );

    \I__7452\ : Span4Mux_v
    port map (
            O => \N__38659\,
            I => \N__38652\
        );

    \I__7451\ : Span4Mux_v
    port map (
            O => \N__38656\,
            I => \N__38649\
        );

    \I__7450\ : InMux
    port map (
            O => \N__38655\,
            I => \N__38646\
        );

    \I__7449\ : Odrv4
    port map (
            O => \N__38652\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__7448\ : Odrv4
    port map (
            O => \N__38649\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__38646\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__7446\ : InMux
    port map (
            O => \N__38639\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__7445\ : InMux
    port map (
            O => \N__38636\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__7444\ : CascadeMux
    port map (
            O => \N__38633\,
            I => \N__38630\
        );

    \I__7443\ : InMux
    port map (
            O => \N__38630\,
            I => \N__38626\
        );

    \I__7442\ : InMux
    port map (
            O => \N__38629\,
            I => \N__38622\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__38626\,
            I => \N__38619\
        );

    \I__7440\ : InMux
    port map (
            O => \N__38625\,
            I => \N__38616\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__38622\,
            I => \N__38613\
        );

    \I__7438\ : Sp12to4
    port map (
            O => \N__38619\,
            I => \N__38608\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__38616\,
            I => \N__38608\
        );

    \I__7436\ : Span4Mux_v
    port map (
            O => \N__38613\,
            I => \N__38605\
        );

    \I__7435\ : Span12Mux_v
    port map (
            O => \N__38608\,
            I => \N__38601\
        );

    \I__7434\ : Span4Mux_v
    port map (
            O => \N__38605\,
            I => \N__38598\
        );

    \I__7433\ : InMux
    port map (
            O => \N__38604\,
            I => \N__38595\
        );

    \I__7432\ : Odrv12
    port map (
            O => \N__38601\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__7431\ : Odrv4
    port map (
            O => \N__38598\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__38595\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__7429\ : InMux
    port map (
            O => \N__38588\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__7428\ : InMux
    port map (
            O => \N__38585\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__7427\ : InMux
    port map (
            O => \N__38582\,
            I => \N__38578\
        );

    \I__7426\ : InMux
    port map (
            O => \N__38581\,
            I => \N__38575\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__38578\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__38575\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__7423\ : InMux
    port map (
            O => \N__38570\,
            I => \N__38566\
        );

    \I__7422\ : InMux
    port map (
            O => \N__38569\,
            I => \N__38563\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__38566\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__38563\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__7419\ : InMux
    port map (
            O => \N__38558\,
            I => \N__38555\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__38555\,
            I => \N__38552\
        );

    \I__7417\ : Span4Mux_v
    port map (
            O => \N__38552\,
            I => \N__38548\
        );

    \I__7416\ : InMux
    port map (
            O => \N__38551\,
            I => \N__38545\
        );

    \I__7415\ : Span4Mux_h
    port map (
            O => \N__38548\,
            I => \N__38542\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__38545\,
            I => \N__38539\
        );

    \I__7413\ : Span4Mux_h
    port map (
            O => \N__38542\,
            I => \N__38534\
        );

    \I__7412\ : Span4Mux_v
    port map (
            O => \N__38539\,
            I => \N__38534\
        );

    \I__7411\ : Span4Mux_v
    port map (
            O => \N__38534\,
            I => \N__38529\
        );

    \I__7410\ : InMux
    port map (
            O => \N__38533\,
            I => \N__38526\
        );

    \I__7409\ : InMux
    port map (
            O => \N__38532\,
            I => \N__38523\
        );

    \I__7408\ : Span4Mux_v
    port map (
            O => \N__38529\,
            I => \N__38520\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__38526\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__38523\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__7405\ : Odrv4
    port map (
            O => \N__38520\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__7404\ : InMux
    port map (
            O => \N__38513\,
            I => \N__38509\
        );

    \I__7403\ : InMux
    port map (
            O => \N__38512\,
            I => \N__38506\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__38509\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__38506\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__7400\ : InMux
    port map (
            O => \N__38501\,
            I => \N__38498\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__38498\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__7398\ : CascadeMux
    port map (
            O => \N__38495\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24_cascade_\
        );

    \I__7397\ : InMux
    port map (
            O => \N__38492\,
            I => \N__38489\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__38489\,
            I => \N__38486\
        );

    \I__7395\ : Span4Mux_h
    port map (
            O => \N__38486\,
            I => \N__38483\
        );

    \I__7394\ : Odrv4
    port map (
            O => \N__38483\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24\
        );

    \I__7393\ : InMux
    port map (
            O => \N__38480\,
            I => \N__38476\
        );

    \I__7392\ : InMux
    port map (
            O => \N__38479\,
            I => \N__38473\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__38476\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__38473\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__7389\ : InMux
    port map (
            O => \N__38468\,
            I => \N__38465\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__38465\,
            I => \N__38462\
        );

    \I__7387\ : Span4Mux_h
    port map (
            O => \N__38462\,
            I => \N__38459\
        );

    \I__7386\ : Odrv4
    port map (
            O => \N__38459\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27\
        );

    \I__7385\ : InMux
    port map (
            O => \N__38456\,
            I => \N__38452\
        );

    \I__7384\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38449\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__38452\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__38449\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__7381\ : CascadeMux
    port map (
            O => \N__38444\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4_cascade_\
        );

    \I__7380\ : InMux
    port map (
            O => \N__38441\,
            I => \N__38438\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__38438\,
            I => \N__38435\
        );

    \I__7378\ : Span4Mux_h
    port map (
            O => \N__38435\,
            I => \N__38432\
        );

    \I__7377\ : Odrv4
    port map (
            O => \N__38432\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4\
        );

    \I__7376\ : InMux
    port map (
            O => \N__38429\,
            I => \N__38426\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__38426\,
            I => \N__38422\
        );

    \I__7374\ : InMux
    port map (
            O => \N__38425\,
            I => \N__38419\
        );

    \I__7373\ : Span4Mux_v
    port map (
            O => \N__38422\,
            I => \N__38416\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__38419\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__7371\ : Odrv4
    port map (
            O => \N__38416\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__7370\ : CascadeMux
    port map (
            O => \N__38411\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27_cascade_\
        );

    \I__7369\ : InMux
    port map (
            O => \N__38408\,
            I => \N__38405\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__38405\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\
        );

    \I__7367\ : CascadeMux
    port map (
            O => \N__38402\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\
        );

    \I__7366\ : InMux
    port map (
            O => \N__38399\,
            I => \N__38395\
        );

    \I__7365\ : InMux
    port map (
            O => \N__38398\,
            I => \N__38392\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__38395\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__38392\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__7362\ : InMux
    port map (
            O => \N__38387\,
            I => \N__38383\
        );

    \I__7361\ : InMux
    port map (
            O => \N__38386\,
            I => \N__38380\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__38383\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__38380\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__7358\ : InMux
    port map (
            O => \N__38375\,
            I => \N__38372\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__38372\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__7356\ : CascadeMux
    port map (
            O => \N__38369\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\
        );

    \I__7355\ : InMux
    port map (
            O => \N__38366\,
            I => \N__38363\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__38363\,
            I => \N__38360\
        );

    \I__7353\ : Span4Mux_h
    port map (
            O => \N__38360\,
            I => \N__38357\
        );

    \I__7352\ : Odrv4
    port map (
            O => \N__38357\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14\
        );

    \I__7351\ : InMux
    port map (
            O => \N__38354\,
            I => \N__38350\
        );

    \I__7350\ : InMux
    port map (
            O => \N__38353\,
            I => \N__38347\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__38350\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__38347\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__7347\ : InMux
    port map (
            O => \N__38342\,
            I => \N__38338\
        );

    \I__7346\ : CascadeMux
    port map (
            O => \N__38341\,
            I => \N__38335\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__38338\,
            I => \N__38331\
        );

    \I__7344\ : InMux
    port map (
            O => \N__38335\,
            I => \N__38326\
        );

    \I__7343\ : InMux
    port map (
            O => \N__38334\,
            I => \N__38326\
        );

    \I__7342\ : Span4Mux_v
    port map (
            O => \N__38331\,
            I => \N__38323\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__38326\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__7340\ : Odrv4
    port map (
            O => \N__38323\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__7339\ : InMux
    port map (
            O => \N__38318\,
            I => \N__38314\
        );

    \I__7338\ : InMux
    port map (
            O => \N__38317\,
            I => \N__38311\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__38314\,
            I => \N__38307\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__38311\,
            I => \N__38304\
        );

    \I__7335\ : InMux
    port map (
            O => \N__38310\,
            I => \N__38301\
        );

    \I__7334\ : Span4Mux_v
    port map (
            O => \N__38307\,
            I => \N__38298\
        );

    \I__7333\ : Sp12to4
    port map (
            O => \N__38304\,
            I => \N__38293\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__38301\,
            I => \N__38293\
        );

    \I__7331\ : Odrv4
    port map (
            O => \N__38298\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__7330\ : Odrv12
    port map (
            O => \N__38293\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__7329\ : ClkMux
    port map (
            O => \N__38288\,
            I => \N__38282\
        );

    \I__7328\ : ClkMux
    port map (
            O => \N__38287\,
            I => \N__38282\
        );

    \I__7327\ : GlobalMux
    port map (
            O => \N__38282\,
            I => \N__38279\
        );

    \I__7326\ : gio2CtrlBuf
    port map (
            O => \N__38279\,
            I => delay_hc_input_c_g
        );

    \I__7325\ : InMux
    port map (
            O => \N__38276\,
            I => \N__38273\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__38273\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__7323\ : InMux
    port map (
            O => \N__38270\,
            I => \N__38266\
        );

    \I__7322\ : InMux
    port map (
            O => \N__38269\,
            I => \N__38263\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__38266\,
            I => \N__38259\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__38263\,
            I => \N__38256\
        );

    \I__7319\ : InMux
    port map (
            O => \N__38262\,
            I => \N__38253\
        );

    \I__7318\ : Span4Mux_v
    port map (
            O => \N__38259\,
            I => \N__38248\
        );

    \I__7317\ : Span4Mux_v
    port map (
            O => \N__38256\,
            I => \N__38248\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__38253\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__7315\ : Odrv4
    port map (
            O => \N__38248\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__7314\ : CascadeMux
    port map (
            O => \N__38243\,
            I => \N__38239\
        );

    \I__7313\ : InMux
    port map (
            O => \N__38242\,
            I => \N__38233\
        );

    \I__7312\ : InMux
    port map (
            O => \N__38239\,
            I => \N__38233\
        );

    \I__7311\ : InMux
    port map (
            O => \N__38238\,
            I => \N__38230\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__38233\,
            I => \N__38227\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__38230\,
            I => \N__38224\
        );

    \I__7308\ : Odrv4
    port map (
            O => \N__38227\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__7307\ : Odrv12
    port map (
            O => \N__38224\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__7306\ : InMux
    port map (
            O => \N__38219\,
            I => \N__38216\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__38216\,
            I => \N__38211\
        );

    \I__7304\ : InMux
    port map (
            O => \N__38215\,
            I => \N__38208\
        );

    \I__7303\ : InMux
    port map (
            O => \N__38214\,
            I => \N__38205\
        );

    \I__7302\ : Sp12to4
    port map (
            O => \N__38211\,
            I => \N__38200\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__38208\,
            I => \N__38200\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__38205\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__7299\ : Odrv12
    port map (
            O => \N__38200\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__7298\ : CascadeMux
    port map (
            O => \N__38195\,
            I => \N__38190\
        );

    \I__7297\ : InMux
    port map (
            O => \N__38194\,
            I => \N__38187\
        );

    \I__7296\ : InMux
    port map (
            O => \N__38193\,
            I => \N__38182\
        );

    \I__7295\ : InMux
    port map (
            O => \N__38190\,
            I => \N__38182\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__38187\,
            I => \N__38179\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__38182\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__7292\ : Odrv12
    port map (
            O => \N__38179\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__7291\ : InMux
    port map (
            O => \N__38174\,
            I => \N__38169\
        );

    \I__7290\ : InMux
    port map (
            O => \N__38173\,
            I => \N__38166\
        );

    \I__7289\ : InMux
    port map (
            O => \N__38172\,
            I => \N__38163\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__38169\,
            I => \N__38160\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__38166\,
            I => \N__38157\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__38163\,
            I => \N__38154\
        );

    \I__7285\ : Odrv4
    port map (
            O => \N__38160\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__7284\ : Odrv4
    port map (
            O => \N__38157\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__7283\ : Odrv4
    port map (
            O => \N__38154\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__7282\ : InMux
    port map (
            O => \N__38147\,
            I => \N__38141\
        );

    \I__7281\ : InMux
    port map (
            O => \N__38146\,
            I => \N__38141\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__38141\,
            I => \N__38137\
        );

    \I__7279\ : InMux
    port map (
            O => \N__38140\,
            I => \N__38134\
        );

    \I__7278\ : Sp12to4
    port map (
            O => \N__38137\,
            I => \N__38129\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__38134\,
            I => \N__38129\
        );

    \I__7276\ : Odrv12
    port map (
            O => \N__38129\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__7275\ : CascadeMux
    port map (
            O => \N__38126\,
            I => \N__38121\
        );

    \I__7274\ : InMux
    port map (
            O => \N__38125\,
            I => \N__38117\
        );

    \I__7273\ : InMux
    port map (
            O => \N__38124\,
            I => \N__38114\
        );

    \I__7272\ : InMux
    port map (
            O => \N__38121\,
            I => \N__38111\
        );

    \I__7271\ : InMux
    port map (
            O => \N__38120\,
            I => \N__38108\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__38117\,
            I => \N__38105\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__38114\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__38111\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__38108\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__7266\ : Odrv4
    port map (
            O => \N__38105\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__38096\,
            I => \N__38093\
        );

    \I__7264\ : InMux
    port map (
            O => \N__38093\,
            I => \N__38088\
        );

    \I__7263\ : InMux
    port map (
            O => \N__38092\,
            I => \N__38085\
        );

    \I__7262\ : InMux
    port map (
            O => \N__38091\,
            I => \N__38082\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__38088\,
            I => \N__38075\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__38085\,
            I => \N__38075\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__38082\,
            I => \N__38075\
        );

    \I__7258\ : Odrv12
    port map (
            O => \N__38075\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__7257\ : InMux
    port map (
            O => \N__38072\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__7256\ : InMux
    port map (
            O => \N__38069\,
            I => \bfn_14_16_0_\
        );

    \I__7255\ : InMux
    port map (
            O => \N__38066\,
            I => \N__38063\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__38063\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__7253\ : InMux
    port map (
            O => \N__38060\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__7252\ : InMux
    port map (
            O => \N__38057\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__7251\ : InMux
    port map (
            O => \N__38054\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__7250\ : InMux
    port map (
            O => \N__38051\,
            I => \N__38048\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__38048\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__7248\ : InMux
    port map (
            O => \N__38045\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__7247\ : InMux
    port map (
            O => \N__38042\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__7246\ : InMux
    port map (
            O => \N__38039\,
            I => \N__38034\
        );

    \I__7245\ : InMux
    port map (
            O => \N__38038\,
            I => \N__38031\
        );

    \I__7244\ : InMux
    port map (
            O => \N__38037\,
            I => \N__38028\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__38034\,
            I => \N__38023\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__38031\,
            I => \N__38023\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__38028\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__7240\ : Odrv4
    port map (
            O => \N__38023\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__7239\ : InMux
    port map (
            O => \N__38018\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__7238\ : InMux
    port map (
            O => \N__38015\,
            I => \N__38012\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__38012\,
            I => \N__38009\
        );

    \I__7236\ : Odrv12
    port map (
            O => \N__38009\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__7235\ : InMux
    port map (
            O => \N__38006\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__7234\ : InMux
    port map (
            O => \N__38003\,
            I => \bfn_14_15_0_\
        );

    \I__7233\ : CascadeMux
    port map (
            O => \N__38000\,
            I => \N__37996\
        );

    \I__7232\ : InMux
    port map (
            O => \N__37999\,
            I => \N__37988\
        );

    \I__7231\ : InMux
    port map (
            O => \N__37996\,
            I => \N__37988\
        );

    \I__7230\ : InMux
    port map (
            O => \N__37995\,
            I => \N__37988\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__37988\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__7228\ : InMux
    port map (
            O => \N__37985\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__7227\ : InMux
    port map (
            O => \N__37982\,
            I => \N__37979\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__37979\,
            I => \N__37976\
        );

    \I__7225\ : Span4Mux_v
    port map (
            O => \N__37976\,
            I => \N__37973\
        );

    \I__7224\ : Odrv4
    port map (
            O => \N__37973\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__7223\ : InMux
    port map (
            O => \N__37970\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__7222\ : InMux
    port map (
            O => \N__37967\,
            I => \N__37964\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__37964\,
            I => \N__37961\
        );

    \I__7220\ : Odrv12
    port map (
            O => \N__37961\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__7219\ : InMux
    port map (
            O => \N__37958\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__7218\ : InMux
    port map (
            O => \N__37955\,
            I => \N__37952\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__37952\,
            I => \N__37949\
        );

    \I__7216\ : Odrv4
    port map (
            O => \N__37949\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__7215\ : InMux
    port map (
            O => \N__37946\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__7214\ : InMux
    port map (
            O => \N__37943\,
            I => \N__37940\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__37940\,
            I => \N__37937\
        );

    \I__7212\ : Odrv4
    port map (
            O => \N__37937\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__7211\ : InMux
    port map (
            O => \N__37934\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__7210\ : InMux
    port map (
            O => \N__37931\,
            I => \N__37928\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__37928\,
            I => \N__37925\
        );

    \I__7208\ : Odrv4
    port map (
            O => \N__37925\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__7207\ : InMux
    port map (
            O => \N__37922\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__7206\ : InMux
    port map (
            O => \N__37919\,
            I => \N__37916\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__37916\,
            I => \N__37913\
        );

    \I__7204\ : Odrv4
    port map (
            O => \N__37913\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__7203\ : InMux
    port map (
            O => \N__37910\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__7202\ : InMux
    port map (
            O => \N__37907\,
            I => \N__37904\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__37904\,
            I => \N__37901\
        );

    \I__7200\ : Odrv4
    port map (
            O => \N__37901\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__7199\ : InMux
    port map (
            O => \N__37898\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__7198\ : InMux
    port map (
            O => \N__37895\,
            I => \bfn_14_14_0_\
        );

    \I__7197\ : InMux
    port map (
            O => \N__37892\,
            I => \N__37889\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__37889\,
            I => \N__37886\
        );

    \I__7195\ : Odrv12
    port map (
            O => \N__37886\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__7194\ : InMux
    port map (
            O => \N__37883\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__7193\ : InMux
    port map (
            O => \N__37880\,
            I => \N__37877\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__37877\,
            I => \N__37874\
        );

    \I__7191\ : Odrv4
    port map (
            O => \N__37874\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__7190\ : InMux
    port map (
            O => \N__37871\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__7189\ : InMux
    port map (
            O => \N__37868\,
            I => \N__37865\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__37865\,
            I => \N__37862\
        );

    \I__7187\ : Odrv4
    port map (
            O => \N__37862\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__7186\ : InMux
    port map (
            O => \N__37859\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__7185\ : InMux
    port map (
            O => \N__37856\,
            I => \N__37853\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__37853\,
            I => \N__37850\
        );

    \I__7183\ : Span4Mux_v
    port map (
            O => \N__37850\,
            I => \N__37847\
        );

    \I__7182\ : Odrv4
    port map (
            O => \N__37847\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__7181\ : InMux
    port map (
            O => \N__37844\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__7180\ : InMux
    port map (
            O => \N__37841\,
            I => \N__37838\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__37838\,
            I => \N__37835\
        );

    \I__7178\ : Odrv12
    port map (
            O => \N__37835\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__7177\ : InMux
    port map (
            O => \N__37832\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__7176\ : InMux
    port map (
            O => \N__37829\,
            I => \N__37826\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__37826\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__7174\ : CascadeMux
    port map (
            O => \N__37823\,
            I => \N__37817\
        );

    \I__7173\ : InMux
    port map (
            O => \N__37822\,
            I => \N__37814\
        );

    \I__7172\ : InMux
    port map (
            O => \N__37821\,
            I => \N__37811\
        );

    \I__7171\ : InMux
    port map (
            O => \N__37820\,
            I => \N__37808\
        );

    \I__7170\ : InMux
    port map (
            O => \N__37817\,
            I => \N__37805\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__37814\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__37811\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__37808\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__37805\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__7165\ : InMux
    port map (
            O => \N__37796\,
            I => \N__37793\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__37793\,
            I => \N__37790\
        );

    \I__7163\ : Odrv4
    port map (
            O => \N__37790\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__7162\ : InMux
    port map (
            O => \N__37787\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__7161\ : InMux
    port map (
            O => \N__37784\,
            I => \N__37781\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__37781\,
            I => \N__37778\
        );

    \I__7159\ : Odrv4
    port map (
            O => \N__37778\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__7158\ : InMux
    port map (
            O => \N__37775\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__7157\ : InMux
    port map (
            O => \N__37772\,
            I => \N__37769\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__37769\,
            I => \N__37766\
        );

    \I__7155\ : Odrv4
    port map (
            O => \N__37766\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__7154\ : InMux
    port map (
            O => \N__37763\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__7153\ : InMux
    port map (
            O => \N__37760\,
            I => \N__37757\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__37757\,
            I => \N__37754\
        );

    \I__7151\ : Odrv4
    port map (
            O => \N__37754\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__7150\ : InMux
    port map (
            O => \N__37751\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__7149\ : InMux
    port map (
            O => \N__37748\,
            I => \N__37745\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__37745\,
            I => \N__37742\
        );

    \I__7147\ : Odrv4
    port map (
            O => \N__37742\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__7146\ : InMux
    port map (
            O => \N__37739\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__7145\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37732\
        );

    \I__7144\ : InMux
    port map (
            O => \N__37735\,
            I => \N__37726\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__37732\,
            I => \N__37723\
        );

    \I__7142\ : InMux
    port map (
            O => \N__37731\,
            I => \N__37720\
        );

    \I__7141\ : CascadeMux
    port map (
            O => \N__37730\,
            I => \N__37716\
        );

    \I__7140\ : InMux
    port map (
            O => \N__37729\,
            I => \N__37713\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__37726\,
            I => \N__37710\
        );

    \I__7138\ : Span4Mux_v
    port map (
            O => \N__37723\,
            I => \N__37707\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__37720\,
            I => \N__37704\
        );

    \I__7136\ : InMux
    port map (
            O => \N__37719\,
            I => \N__37701\
        );

    \I__7135\ : InMux
    port map (
            O => \N__37716\,
            I => \N__37698\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__37713\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__7133\ : Odrv4
    port map (
            O => \N__37710\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__7132\ : Odrv4
    port map (
            O => \N__37707\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__7131\ : Odrv12
    port map (
            O => \N__37704\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__37701\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__37698\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__7128\ : InMux
    port map (
            O => \N__37685\,
            I => \N__37682\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__37682\,
            I => \N__37677\
        );

    \I__7126\ : CascadeMux
    port map (
            O => \N__37681\,
            I => \N__37674\
        );

    \I__7125\ : InMux
    port map (
            O => \N__37680\,
            I => \N__37671\
        );

    \I__7124\ : Span4Mux_v
    port map (
            O => \N__37677\,
            I => \N__37668\
        );

    \I__7123\ : InMux
    port map (
            O => \N__37674\,
            I => \N__37665\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__37671\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\
        );

    \I__7121\ : Odrv4
    port map (
            O => \N__37668\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__37665\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\
        );

    \I__7119\ : InMux
    port map (
            O => \N__37658\,
            I => \N__37655\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__37655\,
            I => \N__37652\
        );

    \I__7117\ : Odrv12
    port map (
            O => \N__37652\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_0\
        );

    \I__7116\ : CEMux
    port map (
            O => \N__37649\,
            I => \N__37644\
        );

    \I__7115\ : CEMux
    port map (
            O => \N__37648\,
            I => \N__37639\
        );

    \I__7114\ : CEMux
    port map (
            O => \N__37647\,
            I => \N__37636\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__37644\,
            I => \N__37632\
        );

    \I__7112\ : CEMux
    port map (
            O => \N__37643\,
            I => \N__37629\
        );

    \I__7111\ : CEMux
    port map (
            O => \N__37642\,
            I => \N__37626\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__37639\,
            I => \N__37623\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__37636\,
            I => \N__37619\
        );

    \I__7108\ : CEMux
    port map (
            O => \N__37635\,
            I => \N__37616\
        );

    \I__7107\ : Span4Mux_h
    port map (
            O => \N__37632\,
            I => \N__37613\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__37629\,
            I => \N__37610\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__37626\,
            I => \N__37607\
        );

    \I__7104\ : Span4Mux_h
    port map (
            O => \N__37623\,
            I => \N__37604\
        );

    \I__7103\ : CEMux
    port map (
            O => \N__37622\,
            I => \N__37601\
        );

    \I__7102\ : Span4Mux_v
    port map (
            O => \N__37619\,
            I => \N__37595\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__37616\,
            I => \N__37595\
        );

    \I__7100\ : Span4Mux_v
    port map (
            O => \N__37613\,
            I => \N__37590\
        );

    \I__7099\ : Span4Mux_h
    port map (
            O => \N__37610\,
            I => \N__37590\
        );

    \I__7098\ : Span4Mux_v
    port map (
            O => \N__37607\,
            I => \N__37587\
        );

    \I__7097\ : Sp12to4
    port map (
            O => \N__37604\,
            I => \N__37582\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__37601\,
            I => \N__37582\
        );

    \I__7095\ : CEMux
    port map (
            O => \N__37600\,
            I => \N__37579\
        );

    \I__7094\ : Odrv4
    port map (
            O => \N__37595\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__7093\ : Odrv4
    port map (
            O => \N__37590\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__7092\ : Odrv4
    port map (
            O => \N__37587\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__7091\ : Odrv12
    port map (
            O => \N__37582\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__37579\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__7089\ : CascadeMux
    port map (
            O => \N__37568\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\
        );

    \I__7088\ : InMux
    port map (
            O => \N__37565\,
            I => \N__37562\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__37562\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17\
        );

    \I__7086\ : InMux
    port map (
            O => \N__37559\,
            I => \N__37556\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__37556\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18\
        );

    \I__7084\ : InMux
    port map (
            O => \N__37553\,
            I => \N__37550\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__37550\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25\
        );

    \I__7082\ : CascadeMux
    port map (
            O => \N__37547\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\
        );

    \I__7081\ : InMux
    port map (
            O => \N__37544\,
            I => \N__37541\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__37541\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9\
        );

    \I__7079\ : InMux
    port map (
            O => \N__37538\,
            I => \N__37535\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__37535\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__37532\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\
        );

    \I__7076\ : InMux
    port map (
            O => \N__37529\,
            I => \N__37526\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__37526\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23\
        );

    \I__7074\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37520\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__37520\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28\
        );

    \I__7072\ : InMux
    port map (
            O => \N__37517\,
            I => \N__37514\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__37514\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__7070\ : CascadeMux
    port map (
            O => \N__37511\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21_cascade_\
        );

    \I__7069\ : InMux
    port map (
            O => \N__37508\,
            I => \N__37505\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__37505\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21\
        );

    \I__7067\ : InMux
    port map (
            O => \N__37502\,
            I => \N__37499\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__37499\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29\
        );

    \I__7065\ : InMux
    port map (
            O => \N__37496\,
            I => \N__37493\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__37493\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__7063\ : InMux
    port map (
            O => \N__37490\,
            I => \N__37487\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__37487\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13\
        );

    \I__7061\ : InMux
    port map (
            O => \N__37484\,
            I => \N__37480\
        );

    \I__7060\ : InMux
    port map (
            O => \N__37483\,
            I => \N__37477\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__37480\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__37477\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__7057\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37468\
        );

    \I__7056\ : InMux
    port map (
            O => \N__37471\,
            I => \N__37465\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__37468\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__37465\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__7053\ : InMux
    port map (
            O => \N__37460\,
            I => \N__37457\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__37457\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__7051\ : CascadeMux
    port map (
            O => \N__37454\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26_cascade_\
        );

    \I__7050\ : CascadeMux
    port map (
            O => \N__37451\,
            I => \N__37448\
        );

    \I__7049\ : InMux
    port map (
            O => \N__37448\,
            I => \N__37445\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__37445\,
            I => \N__37442\
        );

    \I__7047\ : Odrv4
    port map (
            O => \N__37442\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26\
        );

    \I__7046\ : InMux
    port map (
            O => \N__37439\,
            I => \N__37435\
        );

    \I__7045\ : InMux
    port map (
            O => \N__37438\,
            I => \N__37432\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__37435\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__37432\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__7042\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37424\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__37424\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20\
        );

    \I__7040\ : InMux
    port map (
            O => \N__37421\,
            I => \N__37418\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__37418\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12\
        );

    \I__7038\ : InMux
    port map (
            O => \N__37415\,
            I => \N__37412\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__37412\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19\
        );

    \I__7036\ : InMux
    port map (
            O => \N__37409\,
            I => \N__37406\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__37406\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__7034\ : InMux
    port map (
            O => \N__37403\,
            I => \N__37400\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__37400\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__7032\ : CascadeMux
    port map (
            O => \N__37397\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11_cascade_\
        );

    \I__7031\ : CascadeMux
    port map (
            O => \N__37394\,
            I => \N__37391\
        );

    \I__7030\ : InMux
    port map (
            O => \N__37391\,
            I => \N__37388\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__37388\,
            I => \N__37385\
        );

    \I__7028\ : Odrv4
    port map (
            O => \N__37385\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11\
        );

    \I__7027\ : InMux
    port map (
            O => \N__37382\,
            I => \N__37379\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__37379\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__7025\ : CascadeMux
    port map (
            O => \N__37376\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\
        );

    \I__7024\ : InMux
    port map (
            O => \N__37373\,
            I => \N__37370\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__37370\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7\
        );

    \I__7022\ : InMux
    port map (
            O => \N__37367\,
            I => \N__37364\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__37364\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__7020\ : CascadeMux
    port map (
            O => \N__37361\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\
        );

    \I__7019\ : InMux
    port map (
            O => \N__37358\,
            I => \N__37355\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__37355\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8\
        );

    \I__7017\ : InMux
    port map (
            O => \N__37352\,
            I => \N__37348\
        );

    \I__7016\ : InMux
    port map (
            O => \N__37351\,
            I => \N__37345\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__37348\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__37345\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__7013\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37337\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__37337\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3\
        );

    \I__7011\ : InMux
    port map (
            O => \N__37334\,
            I => \N__37331\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__37331\,
            I => \N__37328\
        );

    \I__7009\ : Span12Mux_s6_h
    port map (
            O => \N__37328\,
            I => \N__37325\
        );

    \I__7008\ : Odrv12
    port map (
            O => \N__37325\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0\
        );

    \I__7007\ : InMux
    port map (
            O => \N__37322\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__7006\ : InMux
    port map (
            O => \N__37319\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__7005\ : InMux
    port map (
            O => \N__37316\,
            I => \N__37313\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__37313\,
            I => \N__37310\
        );

    \I__7003\ : Span12Mux_s5_h
    port map (
            O => \N__37310\,
            I => \N__37307\
        );

    \I__7002\ : Odrv12
    port map (
            O => \N__37307\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_CO\
        );

    \I__7001\ : InMux
    port map (
            O => \N__37304\,
            I => \N__37301\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__37301\,
            I => \N__37297\
        );

    \I__6999\ : InMux
    port map (
            O => \N__37300\,
            I => \N__37294\
        );

    \I__6998\ : Span4Mux_v
    port map (
            O => \N__37297\,
            I => \N__37288\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__37294\,
            I => \N__37288\
        );

    \I__6996\ : InMux
    port map (
            O => \N__37293\,
            I => \N__37284\
        );

    \I__6995\ : Span4Mux_v
    port map (
            O => \N__37288\,
            I => \N__37281\
        );

    \I__6994\ : CascadeMux
    port map (
            O => \N__37287\,
            I => \N__37278\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__37284\,
            I => \N__37273\
        );

    \I__6992\ : Span4Mux_h
    port map (
            O => \N__37281\,
            I => \N__37270\
        );

    \I__6991\ : InMux
    port map (
            O => \N__37278\,
            I => \N__37263\
        );

    \I__6990\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37263\
        );

    \I__6989\ : InMux
    port map (
            O => \N__37276\,
            I => \N__37263\
        );

    \I__6988\ : Span12Mux_v
    port map (
            O => \N__37273\,
            I => \N__37260\
        );

    \I__6987\ : Span4Mux_v
    port map (
            O => \N__37270\,
            I => \N__37257\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__37263\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6985\ : Odrv12
    port map (
            O => \N__37260\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6984\ : Odrv4
    port map (
            O => \N__37257\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6983\ : InMux
    port map (
            O => \N__37250\,
            I => \N__37244\
        );

    \I__6982\ : InMux
    port map (
            O => \N__37249\,
            I => \N__37244\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__37244\,
            I => \N__37239\
        );

    \I__6980\ : InMux
    port map (
            O => \N__37243\,
            I => \N__37235\
        );

    \I__6979\ : InMux
    port map (
            O => \N__37242\,
            I => \N__37232\
        );

    \I__6978\ : Span12Mux_h
    port map (
            O => \N__37239\,
            I => \N__37228\
        );

    \I__6977\ : InMux
    port map (
            O => \N__37238\,
            I => \N__37225\
        );

    \I__6976\ : LocalMux
    port map (
            O => \N__37235\,
            I => \N__37222\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__37232\,
            I => \N__37219\
        );

    \I__6974\ : InMux
    port map (
            O => \N__37231\,
            I => \N__37216\
        );

    \I__6973\ : Span12Mux_v
    port map (
            O => \N__37228\,
            I => \N__37211\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__37225\,
            I => \N__37211\
        );

    \I__6971\ : Span4Mux_v
    port map (
            O => \N__37222\,
            I => \N__37206\
        );

    \I__6970\ : Span4Mux_v
    port map (
            O => \N__37219\,
            I => \N__37206\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__37216\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6968\ : Odrv12
    port map (
            O => \N__37211\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6967\ : Odrv4
    port map (
            O => \N__37206\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6966\ : InMux
    port map (
            O => \N__37199\,
            I => \N__37195\
        );

    \I__6965\ : InMux
    port map (
            O => \N__37198\,
            I => \N__37192\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__37195\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__37192\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__6962\ : InMux
    port map (
            O => \N__37187\,
            I => \N__37184\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__37184\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__6960\ : CascadeMux
    port map (
            O => \N__37181\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\
        );

    \I__6959\ : InMux
    port map (
            O => \N__37178\,
            I => \N__37175\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__37175\,
            I => \N__37172\
        );

    \I__6957\ : Odrv4
    port map (
            O => \N__37172\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10\
        );

    \I__6956\ : InMux
    port map (
            O => \N__37169\,
            I => \N__37166\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__37166\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6\
        );

    \I__6954\ : InMux
    port map (
            O => \N__37163\,
            I => \N__37160\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__37160\,
            I => \N__37157\
        );

    \I__6952\ : Span4Mux_v
    port map (
            O => \N__37157\,
            I => \N__37154\
        );

    \I__6951\ : Span4Mux_h
    port map (
            O => \N__37154\,
            I => \N__37151\
        );

    \I__6950\ : Span4Mux_h
    port map (
            O => \N__37151\,
            I => \N__37148\
        );

    \I__6949\ : Span4Mux_h
    port map (
            O => \N__37148\,
            I => \N__37145\
        );

    \I__6948\ : Odrv4
    port map (
            O => \N__37145\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__6947\ : InMux
    port map (
            O => \N__37142\,
            I => \N__37139\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__37139\,
            I => \N__37136\
        );

    \I__6945\ : Span12Mux_s5_h
    port map (
            O => \N__37136\,
            I => \N__37133\
        );

    \I__6944\ : Odrv12
    port map (
            O => \N__37133\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0\
        );

    \I__6943\ : InMux
    port map (
            O => \N__37130\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__6942\ : CascadeMux
    port map (
            O => \N__37127\,
            I => \N__37124\
        );

    \I__6941\ : InMux
    port map (
            O => \N__37124\,
            I => \N__37121\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__37121\,
            I => \N__37118\
        );

    \I__6939\ : Span4Mux_v
    port map (
            O => \N__37118\,
            I => \N__37115\
        );

    \I__6938\ : Span4Mux_v
    port map (
            O => \N__37115\,
            I => \N__37112\
        );

    \I__6937\ : Sp12to4
    port map (
            O => \N__37112\,
            I => \N__37109\
        );

    \I__6936\ : Odrv12
    port map (
            O => \N__37109\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__6935\ : InMux
    port map (
            O => \N__37106\,
            I => \N__37103\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__37103\,
            I => \N__37100\
        );

    \I__6933\ : Span12Mux_s4_h
    port map (
            O => \N__37100\,
            I => \N__37097\
        );

    \I__6932\ : Odrv12
    port map (
            O => \N__37097\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0\
        );

    \I__6931\ : InMux
    port map (
            O => \N__37094\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__6930\ : InMux
    port map (
            O => \N__37091\,
            I => \N__37088\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__37088\,
            I => \N__37085\
        );

    \I__6928\ : Span12Mux_h
    port map (
            O => \N__37085\,
            I => \N__37082\
        );

    \I__6927\ : Span12Mux_h
    port map (
            O => \N__37082\,
            I => \N__37079\
        );

    \I__6926\ : Odrv12
    port map (
            O => \N__37079\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__6925\ : InMux
    port map (
            O => \N__37076\,
            I => \N__37073\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__37073\,
            I => \N__37070\
        );

    \I__6923\ : Span12Mux_s3_h
    port map (
            O => \N__37070\,
            I => \N__37067\
        );

    \I__6922\ : Odrv12
    port map (
            O => \N__37067\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0\
        );

    \I__6921\ : InMux
    port map (
            O => \N__37064\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__37061\,
            I => \N__37058\
        );

    \I__6919\ : InMux
    port map (
            O => \N__37058\,
            I => \N__37055\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__37055\,
            I => \N__37052\
        );

    \I__6917\ : Span4Mux_v
    port map (
            O => \N__37052\,
            I => \N__37049\
        );

    \I__6916\ : Span4Mux_h
    port map (
            O => \N__37049\,
            I => \N__37046\
        );

    \I__6915\ : Span4Mux_h
    port map (
            O => \N__37046\,
            I => \N__37043\
        );

    \I__6914\ : Span4Mux_h
    port map (
            O => \N__37043\,
            I => \N__37040\
        );

    \I__6913\ : Odrv4
    port map (
            O => \N__37040\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__6912\ : InMux
    port map (
            O => \N__37037\,
            I => \N__37034\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__37034\,
            I => \N__37031\
        );

    \I__6910\ : Span12Mux_s2_h
    port map (
            O => \N__37031\,
            I => \N__37028\
        );

    \I__6909\ : Odrv12
    port map (
            O => \N__37028\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0\
        );

    \I__6908\ : InMux
    port map (
            O => \N__37025\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__6907\ : CascadeMux
    port map (
            O => \N__37022\,
            I => \N__37019\
        );

    \I__6906\ : InMux
    port map (
            O => \N__37019\,
            I => \N__37016\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__37016\,
            I => \N__37013\
        );

    \I__6904\ : Span4Mux_v
    port map (
            O => \N__37013\,
            I => \N__37010\
        );

    \I__6903\ : Sp12to4
    port map (
            O => \N__37010\,
            I => \N__37007\
        );

    \I__6902\ : Span12Mux_h
    port map (
            O => \N__37007\,
            I => \N__37004\
        );

    \I__6901\ : Odrv12
    port map (
            O => \N__37004\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__6900\ : InMux
    port map (
            O => \N__37001\,
            I => \N__36998\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__36998\,
            I => \N__36995\
        );

    \I__6898\ : Span12Mux_s9_h
    port map (
            O => \N__36995\,
            I => \N__36992\
        );

    \I__6897\ : Odrv12
    port map (
            O => \N__36992\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0\
        );

    \I__6896\ : InMux
    port map (
            O => \N__36989\,
            I => \bfn_13_22_0_\
        );

    \I__6895\ : InMux
    port map (
            O => \N__36986\,
            I => \N__36983\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__36983\,
            I => \N__36980\
        );

    \I__6893\ : Span4Mux_v
    port map (
            O => \N__36980\,
            I => \N__36977\
        );

    \I__6892\ : Sp12to4
    port map (
            O => \N__36977\,
            I => \N__36974\
        );

    \I__6891\ : Span12Mux_h
    port map (
            O => \N__36974\,
            I => \N__36971\
        );

    \I__6890\ : Odrv12
    port map (
            O => \N__36971\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__6889\ : InMux
    port map (
            O => \N__36968\,
            I => \N__36965\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__36965\,
            I => \N__36962\
        );

    \I__6887\ : Span12Mux_s8_h
    port map (
            O => \N__36962\,
            I => \N__36959\
        );

    \I__6886\ : Odrv12
    port map (
            O => \N__36959\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0\
        );

    \I__6885\ : InMux
    port map (
            O => \N__36956\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__6884\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36950\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__36950\,
            I => \N__36947\
        );

    \I__6882\ : Span4Mux_h
    port map (
            O => \N__36947\,
            I => \N__36944\
        );

    \I__6881\ : Span4Mux_h
    port map (
            O => \N__36944\,
            I => \N__36941\
        );

    \I__6880\ : Sp12to4
    port map (
            O => \N__36941\,
            I => \N__36938\
        );

    \I__6879\ : Span12Mux_v
    port map (
            O => \N__36938\,
            I => \N__36935\
        );

    \I__6878\ : Odrv12
    port map (
            O => \N__36935\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__6877\ : InMux
    port map (
            O => \N__36932\,
            I => \N__36929\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__36929\,
            I => \N__36926\
        );

    \I__6875\ : Span12Mux_s7_h
    port map (
            O => \N__36926\,
            I => \N__36923\
        );

    \I__6874\ : Odrv12
    port map (
            O => \N__36923\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0\
        );

    \I__6873\ : InMux
    port map (
            O => \N__36920\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__6872\ : InMux
    port map (
            O => \N__36917\,
            I => \N__36914\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__36914\,
            I => \N__36911\
        );

    \I__6870\ : Span4Mux_v
    port map (
            O => \N__36911\,
            I => \N__36908\
        );

    \I__6869\ : Sp12to4
    port map (
            O => \N__36908\,
            I => \N__36905\
        );

    \I__6868\ : Span12Mux_h
    port map (
            O => \N__36905\,
            I => \N__36902\
        );

    \I__6867\ : Odrv12
    port map (
            O => \N__36902\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__6866\ : CascadeMux
    port map (
            O => \N__36899\,
            I => \N__36893\
        );

    \I__6865\ : CascadeMux
    port map (
            O => \N__36898\,
            I => \N__36890\
        );

    \I__6864\ : CascadeMux
    port map (
            O => \N__36897\,
            I => \N__36887\
        );

    \I__6863\ : CascadeMux
    port map (
            O => \N__36896\,
            I => \N__36881\
        );

    \I__6862\ : InMux
    port map (
            O => \N__36893\,
            I => \N__36878\
        );

    \I__6861\ : InMux
    port map (
            O => \N__36890\,
            I => \N__36871\
        );

    \I__6860\ : InMux
    port map (
            O => \N__36887\,
            I => \N__36871\
        );

    \I__6859\ : InMux
    port map (
            O => \N__36886\,
            I => \N__36871\
        );

    \I__6858\ : CascadeMux
    port map (
            O => \N__36885\,
            I => \N__36867\
        );

    \I__6857\ : CascadeMux
    port map (
            O => \N__36884\,
            I => \N__36863\
        );

    \I__6856\ : InMux
    port map (
            O => \N__36881\,
            I => \N__36860\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__36878\,
            I => \N__36857\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__36871\,
            I => \N__36854\
        );

    \I__6853\ : InMux
    port map (
            O => \N__36870\,
            I => \N__36845\
        );

    \I__6852\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36845\
        );

    \I__6851\ : InMux
    port map (
            O => \N__36866\,
            I => \N__36845\
        );

    \I__6850\ : InMux
    port map (
            O => \N__36863\,
            I => \N__36845\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__36860\,
            I => \N__36842\
        );

    \I__6848\ : Span4Mux_v
    port map (
            O => \N__36857\,
            I => \N__36835\
        );

    \I__6847\ : Span4Mux_v
    port map (
            O => \N__36854\,
            I => \N__36835\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__36845\,
            I => \N__36835\
        );

    \I__6845\ : Span12Mux_s10_v
    port map (
            O => \N__36842\,
            I => \N__36832\
        );

    \I__6844\ : Span4Mux_v
    port map (
            O => \N__36835\,
            I => \N__36829\
        );

    \I__6843\ : Span12Mux_h
    port map (
            O => \N__36832\,
            I => \N__36826\
        );

    \I__6842\ : Span4Mux_h
    port map (
            O => \N__36829\,
            I => \N__36823\
        );

    \I__6841\ : Span12Mux_h
    port map (
            O => \N__36826\,
            I => \N__36820\
        );

    \I__6840\ : Span4Mux_h
    port map (
            O => \N__36823\,
            I => \N__36817\
        );

    \I__6839\ : Odrv12
    port map (
            O => \N__36820\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__6838\ : Odrv4
    port map (
            O => \N__36817\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__6837\ : InMux
    port map (
            O => \N__36812\,
            I => \N__36809\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__36809\,
            I => \N__36806\
        );

    \I__6835\ : Span4Mux_v
    port map (
            O => \N__36806\,
            I => \N__36803\
        );

    \I__6834\ : Span4Mux_h
    port map (
            O => \N__36803\,
            I => \N__36800\
        );

    \I__6833\ : Span4Mux_h
    port map (
            O => \N__36800\,
            I => \N__36797\
        );

    \I__6832\ : Span4Mux_h
    port map (
            O => \N__36797\,
            I => \N__36794\
        );

    \I__6831\ : Odrv4
    port map (
            O => \N__36794\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__6830\ : CascadeMux
    port map (
            O => \N__36791\,
            I => \N__36788\
        );

    \I__6829\ : InMux
    port map (
            O => \N__36788\,
            I => \N__36785\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__36785\,
            I => \N__36782\
        );

    \I__6827\ : Sp12to4
    port map (
            O => \N__36782\,
            I => \N__36779\
        );

    \I__6826\ : Span12Mux_v
    port map (
            O => \N__36779\,
            I => \N__36776\
        );

    \I__6825\ : Odrv12
    port map (
            O => \N__36776\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__6824\ : CascadeMux
    port map (
            O => \N__36773\,
            I => \N__36770\
        );

    \I__6823\ : InMux
    port map (
            O => \N__36770\,
            I => \N__36767\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__36767\,
            I => \N__36764\
        );

    \I__6821\ : Span12Mux_s9_h
    port map (
            O => \N__36764\,
            I => \N__36761\
        );

    \I__6820\ : Odrv12
    port map (
            O => \N__36761\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_8\
        );

    \I__6819\ : InMux
    port map (
            O => \N__36758\,
            I => \N__36755\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__36755\,
            I => \N__36752\
        );

    \I__6817\ : Span4Mux_v
    port map (
            O => \N__36752\,
            I => \N__36749\
        );

    \I__6816\ : Sp12to4
    port map (
            O => \N__36749\,
            I => \N__36746\
        );

    \I__6815\ : Span12Mux_h
    port map (
            O => \N__36746\,
            I => \N__36743\
        );

    \I__6814\ : Odrv12
    port map (
            O => \N__36743\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__6813\ : CascadeMux
    port map (
            O => \N__36740\,
            I => \N__36737\
        );

    \I__6812\ : InMux
    port map (
            O => \N__36737\,
            I => \N__36734\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__36734\,
            I => \N__36731\
        );

    \I__6810\ : Span12Mux_v
    port map (
            O => \N__36731\,
            I => \N__36728\
        );

    \I__6809\ : Span12Mux_h
    port map (
            O => \N__36728\,
            I => \N__36725\
        );

    \I__6808\ : Odrv12
    port map (
            O => \N__36725\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__6807\ : CascadeMux
    port map (
            O => \N__36722\,
            I => \N__36719\
        );

    \I__6806\ : InMux
    port map (
            O => \N__36719\,
            I => \N__36716\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__36716\,
            I => \N__36713\
        );

    \I__6804\ : Span12Mux_s8_h
    port map (
            O => \N__36713\,
            I => \N__36710\
        );

    \I__6803\ : Odrv12
    port map (
            O => \N__36710\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0\
        );

    \I__6802\ : InMux
    port map (
            O => \N__36707\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__6801\ : InMux
    port map (
            O => \N__36704\,
            I => \N__36701\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__36701\,
            I => \N__36698\
        );

    \I__6799\ : Span4Mux_h
    port map (
            O => \N__36698\,
            I => \N__36695\
        );

    \I__6798\ : Span4Mux_h
    port map (
            O => \N__36695\,
            I => \N__36692\
        );

    \I__6797\ : Sp12to4
    port map (
            O => \N__36692\,
            I => \N__36689\
        );

    \I__6796\ : Span12Mux_v
    port map (
            O => \N__36689\,
            I => \N__36686\
        );

    \I__6795\ : Odrv12
    port map (
            O => \N__36686\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__6794\ : CascadeMux
    port map (
            O => \N__36683\,
            I => \N__36680\
        );

    \I__6793\ : InMux
    port map (
            O => \N__36680\,
            I => \N__36677\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__36677\,
            I => \N__36674\
        );

    \I__6791\ : Span12Mux_v
    port map (
            O => \N__36674\,
            I => \N__36671\
        );

    \I__6790\ : Span12Mux_h
    port map (
            O => \N__36671\,
            I => \N__36668\
        );

    \I__6789\ : Odrv12
    port map (
            O => \N__36668\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__6788\ : CascadeMux
    port map (
            O => \N__36665\,
            I => \N__36662\
        );

    \I__6787\ : InMux
    port map (
            O => \N__36662\,
            I => \N__36659\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__36659\,
            I => \N__36656\
        );

    \I__6785\ : Span12Mux_s7_h
    port map (
            O => \N__36656\,
            I => \N__36653\
        );

    \I__6784\ : Odrv12
    port map (
            O => \N__36653\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0\
        );

    \I__6783\ : InMux
    port map (
            O => \N__36650\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__6782\ : InMux
    port map (
            O => \N__36647\,
            I => \N__36644\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__36644\,
            I => \N__36641\
        );

    \I__6780\ : Span4Mux_v
    port map (
            O => \N__36641\,
            I => \N__36638\
        );

    \I__6779\ : Sp12to4
    port map (
            O => \N__36638\,
            I => \N__36635\
        );

    \I__6778\ : Span12Mux_h
    port map (
            O => \N__36635\,
            I => \N__36632\
        );

    \I__6777\ : Odrv12
    port map (
            O => \N__36632\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__6776\ : CascadeMux
    port map (
            O => \N__36629\,
            I => \N__36626\
        );

    \I__6775\ : InMux
    port map (
            O => \N__36626\,
            I => \N__36623\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__36623\,
            I => \N__36620\
        );

    \I__6773\ : Span4Mux_v
    port map (
            O => \N__36620\,
            I => \N__36617\
        );

    \I__6772\ : Span4Mux_h
    port map (
            O => \N__36617\,
            I => \N__36614\
        );

    \I__6771\ : Span4Mux_h
    port map (
            O => \N__36614\,
            I => \N__36611\
        );

    \I__6770\ : Odrv4
    port map (
            O => \N__36611\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__6769\ : CascadeMux
    port map (
            O => \N__36608\,
            I => \N__36605\
        );

    \I__6768\ : InMux
    port map (
            O => \N__36605\,
            I => \N__36602\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__36602\,
            I => \N__36599\
        );

    \I__6766\ : Span12Mux_s6_h
    port map (
            O => \N__36599\,
            I => \N__36596\
        );

    \I__6765\ : Odrv12
    port map (
            O => \N__36596\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0\
        );

    \I__6764\ : InMux
    port map (
            O => \N__36593\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__6763\ : InMux
    port map (
            O => \N__36590\,
            I => \N__36584\
        );

    \I__6762\ : InMux
    port map (
            O => \N__36589\,
            I => \N__36584\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__36584\,
            I => \N__36579\
        );

    \I__6760\ : InMux
    port map (
            O => \N__36583\,
            I => \N__36576\
        );

    \I__6759\ : InMux
    port map (
            O => \N__36582\,
            I => \N__36573\
        );

    \I__6758\ : Odrv4
    port map (
            O => \N__36579\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__36576\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__36573\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6755\ : CascadeMux
    port map (
            O => \N__36566\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__6754\ : InMux
    port map (
            O => \N__36563\,
            I => \N__36560\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__36560\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__6752\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36553\
        );

    \I__6751\ : InMux
    port map (
            O => \N__36556\,
            I => \N__36550\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__36553\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__36550\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0\
        );

    \I__6748\ : InMux
    port map (
            O => \N__36545\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26\
        );

    \I__6747\ : InMux
    port map (
            O => \N__36542\,
            I => \N__36538\
        );

    \I__6746\ : InMux
    port map (
            O => \N__36541\,
            I => \N__36535\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__36538\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__36535\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0\
        );

    \I__6743\ : InMux
    port map (
            O => \N__36530\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27\
        );

    \I__6742\ : InMux
    port map (
            O => \N__36527\,
            I => \N__36523\
        );

    \I__6741\ : InMux
    port map (
            O => \N__36526\,
            I => \N__36520\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__36523\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__36520\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0\
        );

    \I__6738\ : InMux
    port map (
            O => \N__36515\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28\
        );

    \I__6737\ : InMux
    port map (
            O => \N__36512\,
            I => \N__36508\
        );

    \I__6736\ : InMux
    port map (
            O => \N__36511\,
            I => \N__36505\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__36508\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__36505\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0\
        );

    \I__6733\ : InMux
    port map (
            O => \N__36500\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29\
        );

    \I__6732\ : InMux
    port map (
            O => \N__36497\,
            I => \N__36494\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__36494\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO\
        );

    \I__6730\ : InMux
    port map (
            O => \N__36491\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30\
        );

    \I__6729\ : InMux
    port map (
            O => \N__36488\,
            I => \N__36485\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__36485\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30\
        );

    \I__6727\ : InMux
    port map (
            O => \N__36482\,
            I => \N__36479\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__36479\,
            I => \N__36475\
        );

    \I__6725\ : InMux
    port map (
            O => \N__36478\,
            I => \N__36472\
        );

    \I__6724\ : Odrv4
    port map (
            O => \N__36475\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_28
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__36472\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_28
        );

    \I__6722\ : InMux
    port map (
            O => \N__36467\,
            I => \N__36464\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__36464\,
            I => \N__36461\
        );

    \I__6720\ : Span4Mux_h
    port map (
            O => \N__36461\,
            I => \N__36457\
        );

    \I__6719\ : InMux
    port map (
            O => \N__36460\,
            I => \N__36453\
        );

    \I__6718\ : Span4Mux_v
    port map (
            O => \N__36457\,
            I => \N__36450\
        );

    \I__6717\ : InMux
    port map (
            O => \N__36456\,
            I => \N__36447\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__36453\,
            I => \N__36444\
        );

    \I__6715\ : Span4Mux_v
    port map (
            O => \N__36450\,
            I => \N__36441\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__36447\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_31\
        );

    \I__6713\ : Odrv12
    port map (
            O => \N__36444\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_31\
        );

    \I__6712\ : Odrv4
    port map (
            O => \N__36441\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_31\
        );

    \I__6711\ : InMux
    port map (
            O => \N__36434\,
            I => \N__36431\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__36431\,
            I => \N__36426\
        );

    \I__6709\ : InMux
    port map (
            O => \N__36430\,
            I => \N__36423\
        );

    \I__6708\ : InMux
    port map (
            O => \N__36429\,
            I => \N__36420\
        );

    \I__6707\ : Span12Mux_v
    port map (
            O => \N__36426\,
            I => \N__36417\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__36423\,
            I => \N__36414\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__36420\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_30\
        );

    \I__6704\ : Odrv12
    port map (
            O => \N__36417\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_30\
        );

    \I__6703\ : Odrv12
    port map (
            O => \N__36414\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_30\
        );

    \I__6702\ : InMux
    port map (
            O => \N__36407\,
            I => \N__36398\
        );

    \I__6701\ : InMux
    port map (
            O => \N__36406\,
            I => \N__36398\
        );

    \I__6700\ : InMux
    port map (
            O => \N__36405\,
            I => \N__36398\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__36398\,
            I => \N__36394\
        );

    \I__6698\ : InMux
    port map (
            O => \N__36397\,
            I => \N__36391\
        );

    \I__6697\ : Span4Mux_v
    port map (
            O => \N__36394\,
            I => \N__36388\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__36391\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28\
        );

    \I__6695\ : Odrv4
    port map (
            O => \N__36388\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28\
        );

    \I__6694\ : CascadeMux
    port map (
            O => \N__36383\,
            I => \N__36380\
        );

    \I__6693\ : InMux
    port map (
            O => \N__36380\,
            I => \N__36377\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__36377\,
            I => \N__36374\
        );

    \I__6691\ : Span4Mux_h
    port map (
            O => \N__36374\,
            I => \N__36371\
        );

    \I__6690\ : Odrv4
    port map (
            O => \N__36371\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt30\
        );

    \I__6689\ : InMux
    port map (
            O => \N__36368\,
            I => \N__36364\
        );

    \I__6688\ : InMux
    port map (
            O => \N__36367\,
            I => \N__36361\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__36364\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__36361\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9\
        );

    \I__6685\ : InMux
    port map (
            O => \N__36356\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18\
        );

    \I__6684\ : InMux
    port map (
            O => \N__36353\,
            I => \N__36349\
        );

    \I__6683\ : InMux
    port map (
            O => \N__36352\,
            I => \N__36346\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__36349\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__36346\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9\
        );

    \I__6680\ : InMux
    port map (
            O => \N__36341\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19\
        );

    \I__6679\ : InMux
    port map (
            O => \N__36338\,
            I => \N__36334\
        );

    \I__6678\ : InMux
    port map (
            O => \N__36337\,
            I => \N__36331\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__36334\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__36331\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0\
        );

    \I__6675\ : InMux
    port map (
            O => \N__36326\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20\
        );

    \I__6674\ : InMux
    port map (
            O => \N__36323\,
            I => \N__36320\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__36320\,
            I => \N__36317\
        );

    \I__6672\ : Odrv4
    port map (
            O => \N__36317\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22\
        );

    \I__6671\ : InMux
    port map (
            O => \N__36314\,
            I => \N__36310\
        );

    \I__6670\ : InMux
    port map (
            O => \N__36313\,
            I => \N__36307\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__36310\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__36307\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0\
        );

    \I__6667\ : InMux
    port map (
            O => \N__36302\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21\
        );

    \I__6666\ : InMux
    port map (
            O => \N__36299\,
            I => \N__36295\
        );

    \I__6665\ : InMux
    port map (
            O => \N__36298\,
            I => \N__36292\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__36295\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__36292\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0\
        );

    \I__6662\ : InMux
    port map (
            O => \N__36287\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22\
        );

    \I__6661\ : InMux
    port map (
            O => \N__36284\,
            I => \N__36280\
        );

    \I__6660\ : InMux
    port map (
            O => \N__36283\,
            I => \N__36277\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__36280\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__36277\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0\
        );

    \I__6657\ : InMux
    port map (
            O => \N__36272\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23\
        );

    \I__6656\ : InMux
    port map (
            O => \N__36269\,
            I => \N__36265\
        );

    \I__6655\ : InMux
    port map (
            O => \N__36268\,
            I => \N__36262\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__36265\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__36262\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0\
        );

    \I__6652\ : InMux
    port map (
            O => \N__36257\,
            I => \bfn_13_10_0_\
        );

    \I__6651\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36250\
        );

    \I__6650\ : InMux
    port map (
            O => \N__36253\,
            I => \N__36247\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__36250\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__36247\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0\
        );

    \I__6647\ : InMux
    port map (
            O => \N__36242\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25\
        );

    \I__6646\ : InMux
    port map (
            O => \N__36239\,
            I => \N__36235\
        );

    \I__6645\ : InMux
    port map (
            O => \N__36238\,
            I => \N__36232\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__36235\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__36232\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3\
        );

    \I__6642\ : InMux
    port map (
            O => \N__36227\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9\
        );

    \I__6641\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36220\
        );

    \I__6640\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36217\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__36220\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__36217\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49\
        );

    \I__6637\ : InMux
    port map (
            O => \N__36212\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10\
        );

    \I__6636\ : InMux
    port map (
            O => \N__36209\,
            I => \N__36205\
        );

    \I__6635\ : InMux
    port map (
            O => \N__36208\,
            I => \N__36202\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__36205\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__36202\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59\
        );

    \I__6632\ : InMux
    port map (
            O => \N__36197\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11\
        );

    \I__6631\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36190\
        );

    \I__6630\ : InMux
    port map (
            O => \N__36193\,
            I => \N__36187\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__36190\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__36187\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69\
        );

    \I__6627\ : InMux
    port map (
            O => \N__36182\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12\
        );

    \I__6626\ : InMux
    port map (
            O => \N__36179\,
            I => \N__36175\
        );

    \I__6625\ : InMux
    port map (
            O => \N__36178\,
            I => \N__36172\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__36175\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__36172\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79\
        );

    \I__6622\ : InMux
    port map (
            O => \N__36167\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13\
        );

    \I__6621\ : InMux
    port map (
            O => \N__36164\,
            I => \N__36161\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__36161\,
            I => \N__36158\
        );

    \I__6619\ : Odrv4
    port map (
            O => \N__36158\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15\
        );

    \I__6618\ : InMux
    port map (
            O => \N__36155\,
            I => \N__36151\
        );

    \I__6617\ : InMux
    port map (
            O => \N__36154\,
            I => \N__36148\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__36151\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__36148\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099\
        );

    \I__6614\ : InMux
    port map (
            O => \N__36143\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14\
        );

    \I__6613\ : InMux
    port map (
            O => \N__36140\,
            I => \N__36136\
        );

    \I__6612\ : InMux
    port map (
            O => \N__36139\,
            I => \N__36133\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__36136\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__36133\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9\
        );

    \I__6609\ : InMux
    port map (
            O => \N__36128\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15\
        );

    \I__6608\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36121\
        );

    \I__6607\ : InMux
    port map (
            O => \N__36124\,
            I => \N__36118\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__36121\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__36118\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9\
        );

    \I__6604\ : InMux
    port map (
            O => \N__36113\,
            I => \bfn_13_9_0_\
        );

    \I__6603\ : InMux
    port map (
            O => \N__36110\,
            I => \N__36106\
        );

    \I__6602\ : InMux
    port map (
            O => \N__36109\,
            I => \N__36103\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__36106\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__36103\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9\
        );

    \I__6599\ : InMux
    port map (
            O => \N__36098\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17\
        );

    \I__6598\ : InMux
    port map (
            O => \N__36095\,
            I => \N__36092\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__36092\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2\
        );

    \I__6596\ : InMux
    port map (
            O => \N__36089\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2\
        );

    \I__6595\ : InMux
    port map (
            O => \N__36086\,
            I => \N__36082\
        );

    \I__6594\ : InMux
    port map (
            O => \N__36085\,
            I => \N__36079\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__36082\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__36079\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0\
        );

    \I__6591\ : InMux
    port map (
            O => \N__36074\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3\
        );

    \I__6590\ : InMux
    port map (
            O => \N__36071\,
            I => \N__36068\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__36068\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5\
        );

    \I__6588\ : InMux
    port map (
            O => \N__36065\,
            I => \N__36061\
        );

    \I__6587\ : InMux
    port map (
            O => \N__36064\,
            I => \N__36058\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__36061\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__36058\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0\
        );

    \I__6584\ : InMux
    port map (
            O => \N__36053\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4\
        );

    \I__6583\ : InMux
    port map (
            O => \N__36050\,
            I => \N__36046\
        );

    \I__6582\ : InMux
    port map (
            O => \N__36049\,
            I => \N__36043\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__36046\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__36043\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0\
        );

    \I__6579\ : InMux
    port map (
            O => \N__36038\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5\
        );

    \I__6578\ : InMux
    port map (
            O => \N__36035\,
            I => \N__36031\
        );

    \I__6577\ : InMux
    port map (
            O => \N__36034\,
            I => \N__36028\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__36031\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__36028\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26\
        );

    \I__6574\ : InMux
    port map (
            O => \N__36023\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6\
        );

    \I__6573\ : InMux
    port map (
            O => \N__36020\,
            I => \N__36016\
        );

    \I__6572\ : InMux
    port map (
            O => \N__36019\,
            I => \N__36013\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__36016\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__36013\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381\
        );

    \I__6569\ : InMux
    port map (
            O => \N__36008\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7\
        );

    \I__6568\ : InMux
    port map (
            O => \N__36005\,
            I => \N__36001\
        );

    \I__6567\ : InMux
    port map (
            O => \N__36004\,
            I => \N__35998\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__36001\,
            I => \N__35993\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__35998\,
            I => \N__35993\
        );

    \I__6564\ : Odrv4
    port map (
            O => \N__35993\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2\
        );

    \I__6563\ : InMux
    port map (
            O => \N__35990\,
            I => \bfn_13_8_0_\
        );

    \I__6562\ : CascadeMux
    port map (
            O => \N__35987\,
            I => \N__35977\
        );

    \I__6561\ : CascadeMux
    port map (
            O => \N__35986\,
            I => \N__35974\
        );

    \I__6560\ : CascadeMux
    port map (
            O => \N__35985\,
            I => \N__35970\
        );

    \I__6559\ : CascadeMux
    port map (
            O => \N__35984\,
            I => \N__35967\
        );

    \I__6558\ : CascadeMux
    port map (
            O => \N__35983\,
            I => \N__35964\
        );

    \I__6557\ : CascadeMux
    port map (
            O => \N__35982\,
            I => \N__35959\
        );

    \I__6556\ : CascadeMux
    port map (
            O => \N__35981\,
            I => \N__35955\
        );

    \I__6555\ : InMux
    port map (
            O => \N__35980\,
            I => \N__35952\
        );

    \I__6554\ : InMux
    port map (
            O => \N__35977\,
            I => \N__35947\
        );

    \I__6553\ : InMux
    port map (
            O => \N__35974\,
            I => \N__35947\
        );

    \I__6552\ : InMux
    port map (
            O => \N__35973\,
            I => \N__35936\
        );

    \I__6551\ : InMux
    port map (
            O => \N__35970\,
            I => \N__35936\
        );

    \I__6550\ : InMux
    port map (
            O => \N__35967\,
            I => \N__35936\
        );

    \I__6549\ : InMux
    port map (
            O => \N__35964\,
            I => \N__35936\
        );

    \I__6548\ : InMux
    port map (
            O => \N__35963\,
            I => \N__35936\
        );

    \I__6547\ : InMux
    port map (
            O => \N__35962\,
            I => \N__35927\
        );

    \I__6546\ : InMux
    port map (
            O => \N__35959\,
            I => \N__35927\
        );

    \I__6545\ : InMux
    port map (
            O => \N__35958\,
            I => \N__35927\
        );

    \I__6544\ : InMux
    port map (
            O => \N__35955\,
            I => \N__35927\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__35952\,
            I => \N__35924\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__35947\,
            I => \N__35917\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__35936\,
            I => \N__35917\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__35927\,
            I => \N__35917\
        );

    \I__6539\ : Span4Mux_v
    port map (
            O => \N__35924\,
            I => \N__35914\
        );

    \I__6538\ : Span4Mux_v
    port map (
            O => \N__35917\,
            I => \N__35911\
        );

    \I__6537\ : Sp12to4
    port map (
            O => \N__35914\,
            I => \N__35906\
        );

    \I__6536\ : Sp12to4
    port map (
            O => \N__35911\,
            I => \N__35906\
        );

    \I__6535\ : Span12Mux_h
    port map (
            O => \N__35906\,
            I => \N__35903\
        );

    \I__6534\ : Odrv12
    port map (
            O => \N__35903\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__6533\ : CascadeMux
    port map (
            O => \N__35900\,
            I => \N__35897\
        );

    \I__6532\ : InMux
    port map (
            O => \N__35897\,
            I => \N__35894\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__35894\,
            I => \N__35891\
        );

    \I__6530\ : Span12Mux_v
    port map (
            O => \N__35891\,
            I => \N__35888\
        );

    \I__6529\ : Span12Mux_h
    port map (
            O => \N__35888\,
            I => \N__35885\
        );

    \I__6528\ : Odrv12
    port map (
            O => \N__35885\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_14\
        );

    \I__6527\ : InMux
    port map (
            O => \N__35882\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\
        );

    \I__6526\ : InMux
    port map (
            O => \N__35879\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\
        );

    \I__6525\ : IoInMux
    port map (
            O => \N__35876\,
            I => \N__35873\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__35873\,
            I => \N__35870\
        );

    \I__6523\ : Span4Mux_s0_v
    port map (
            O => \N__35870\,
            I => \N__35867\
        );

    \I__6522\ : Odrv4
    port map (
            O => \N__35867\,
            I => \GB_BUFFER_red_c_g_THRU_CO\
        );

    \I__6521\ : InMux
    port map (
            O => \N__35864\,
            I => \N__35861\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__35861\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__6519\ : CascadeMux
    port map (
            O => \N__35858\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15_cascade_\
        );

    \I__6518\ : InMux
    port map (
            O => \N__35855\,
            I => \N__35852\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__35852\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1\
        );

    \I__6516\ : CascadeMux
    port map (
            O => \N__35849\,
            I => \N__35846\
        );

    \I__6515\ : InMux
    port map (
            O => \N__35846\,
            I => \N__35843\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__35843\,
            I => \N__35840\
        );

    \I__6513\ : Sp12to4
    port map (
            O => \N__35840\,
            I => \N__35837\
        );

    \I__6512\ : Span12Mux_v
    port map (
            O => \N__35837\,
            I => \N__35834\
        );

    \I__6511\ : Span12Mux_h
    port map (
            O => \N__35834\,
            I => \N__35831\
        );

    \I__6510\ : Odrv12
    port map (
            O => \N__35831\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_5\
        );

    \I__6509\ : InMux
    port map (
            O => \N__35828\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\
        );

    \I__6508\ : InMux
    port map (
            O => \N__35825\,
            I => \N__35822\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__35822\,
            I => \N__35819\
        );

    \I__6506\ : Span12Mux_v
    port map (
            O => \N__35819\,
            I => \N__35816\
        );

    \I__6505\ : Span12Mux_h
    port map (
            O => \N__35816\,
            I => \N__35813\
        );

    \I__6504\ : Odrv12
    port map (
            O => \N__35813\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_6\
        );

    \I__6503\ : InMux
    port map (
            O => \N__35810\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\
        );

    \I__6502\ : CascadeMux
    port map (
            O => \N__35807\,
            I => \N__35804\
        );

    \I__6501\ : InMux
    port map (
            O => \N__35804\,
            I => \N__35801\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__35801\,
            I => \N__35798\
        );

    \I__6499\ : Span4Mux_v
    port map (
            O => \N__35798\,
            I => \N__35795\
        );

    \I__6498\ : Sp12to4
    port map (
            O => \N__35795\,
            I => \N__35792\
        );

    \I__6497\ : Span12Mux_v
    port map (
            O => \N__35792\,
            I => \N__35789\
        );

    \I__6496\ : Span12Mux_h
    port map (
            O => \N__35789\,
            I => \N__35786\
        );

    \I__6495\ : Odrv12
    port map (
            O => \N__35786\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_7\
        );

    \I__6494\ : InMux
    port map (
            O => \N__35783\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\
        );

    \I__6493\ : CascadeMux
    port map (
            O => \N__35780\,
            I => \N__35777\
        );

    \I__6492\ : InMux
    port map (
            O => \N__35777\,
            I => \N__35774\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__35774\,
            I => \N__35771\
        );

    \I__6490\ : Span12Mux_s11_v
    port map (
            O => \N__35771\,
            I => \N__35768\
        );

    \I__6489\ : Span12Mux_h
    port map (
            O => \N__35768\,
            I => \N__35765\
        );

    \I__6488\ : Odrv12
    port map (
            O => \N__35765\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_8\
        );

    \I__6487\ : InMux
    port map (
            O => \N__35762\,
            I => \bfn_12_24_0_\
        );

    \I__6486\ : InMux
    port map (
            O => \N__35759\,
            I => \N__35756\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__35756\,
            I => \N__35753\
        );

    \I__6484\ : Span4Mux_v
    port map (
            O => \N__35753\,
            I => \N__35750\
        );

    \I__6483\ : Sp12to4
    port map (
            O => \N__35750\,
            I => \N__35747\
        );

    \I__6482\ : Span12Mux_h
    port map (
            O => \N__35747\,
            I => \N__35744\
        );

    \I__6481\ : Odrv12
    port map (
            O => \N__35744\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_9\
        );

    \I__6480\ : InMux
    port map (
            O => \N__35741\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\
        );

    \I__6479\ : InMux
    port map (
            O => \N__35738\,
            I => \N__35735\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__35735\,
            I => \N__35732\
        );

    \I__6477\ : Span12Mux_v
    port map (
            O => \N__35732\,
            I => \N__35729\
        );

    \I__6476\ : Span12Mux_h
    port map (
            O => \N__35729\,
            I => \N__35726\
        );

    \I__6475\ : Odrv12
    port map (
            O => \N__35726\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_10\
        );

    \I__6474\ : InMux
    port map (
            O => \N__35723\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\
        );

    \I__6473\ : InMux
    port map (
            O => \N__35720\,
            I => \N__35717\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__35717\,
            I => \N__35714\
        );

    \I__6471\ : Span12Mux_v
    port map (
            O => \N__35714\,
            I => \N__35711\
        );

    \I__6470\ : Span12Mux_h
    port map (
            O => \N__35711\,
            I => \N__35708\
        );

    \I__6469\ : Odrv12
    port map (
            O => \N__35708\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_11\
        );

    \I__6468\ : InMux
    port map (
            O => \N__35705\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\
        );

    \I__6467\ : InMux
    port map (
            O => \N__35702\,
            I => \N__35699\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__35699\,
            I => \N__35696\
        );

    \I__6465\ : Span12Mux_v
    port map (
            O => \N__35696\,
            I => \N__35693\
        );

    \I__6464\ : Span12Mux_h
    port map (
            O => \N__35693\,
            I => \N__35690\
        );

    \I__6463\ : Odrv12
    port map (
            O => \N__35690\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_12\
        );

    \I__6462\ : InMux
    port map (
            O => \N__35687\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\
        );

    \I__6461\ : InMux
    port map (
            O => \N__35684\,
            I => \N__35681\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__35681\,
            I => \N__35678\
        );

    \I__6459\ : Span12Mux_v
    port map (
            O => \N__35678\,
            I => \N__35675\
        );

    \I__6458\ : Span12Mux_h
    port map (
            O => \N__35675\,
            I => \N__35672\
        );

    \I__6457\ : Odrv12
    port map (
            O => \N__35672\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_13\
        );

    \I__6456\ : InMux
    port map (
            O => \N__35669\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__35666\,
            I => \N__35663\
        );

    \I__6454\ : InMux
    port map (
            O => \N__35663\,
            I => \N__35658\
        );

    \I__6453\ : InMux
    port map (
            O => \N__35662\,
            I => \N__35655\
        );

    \I__6452\ : InMux
    port map (
            O => \N__35661\,
            I => \N__35652\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__35658\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__35655\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__35652\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__6448\ : InMux
    port map (
            O => \N__35645\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__35642\,
            I => \N__35638\
        );

    \I__6446\ : InMux
    port map (
            O => \N__35641\,
            I => \N__35635\
        );

    \I__6445\ : InMux
    port map (
            O => \N__35638\,
            I => \N__35632\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__35635\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__35632\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__6442\ : InMux
    port map (
            O => \N__35627\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__6441\ : InMux
    port map (
            O => \N__35624\,
            I => \N__35590\
        );

    \I__6440\ : InMux
    port map (
            O => \N__35623\,
            I => \N__35590\
        );

    \I__6439\ : InMux
    port map (
            O => \N__35622\,
            I => \N__35590\
        );

    \I__6438\ : InMux
    port map (
            O => \N__35621\,
            I => \N__35590\
        );

    \I__6437\ : InMux
    port map (
            O => \N__35620\,
            I => \N__35581\
        );

    \I__6436\ : InMux
    port map (
            O => \N__35619\,
            I => \N__35581\
        );

    \I__6435\ : InMux
    port map (
            O => \N__35618\,
            I => \N__35572\
        );

    \I__6434\ : InMux
    port map (
            O => \N__35617\,
            I => \N__35572\
        );

    \I__6433\ : InMux
    port map (
            O => \N__35616\,
            I => \N__35572\
        );

    \I__6432\ : InMux
    port map (
            O => \N__35615\,
            I => \N__35572\
        );

    \I__6431\ : InMux
    port map (
            O => \N__35614\,
            I => \N__35563\
        );

    \I__6430\ : InMux
    port map (
            O => \N__35613\,
            I => \N__35563\
        );

    \I__6429\ : InMux
    port map (
            O => \N__35612\,
            I => \N__35563\
        );

    \I__6428\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35563\
        );

    \I__6427\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35554\
        );

    \I__6426\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35554\
        );

    \I__6425\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35554\
        );

    \I__6424\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35554\
        );

    \I__6423\ : InMux
    port map (
            O => \N__35606\,
            I => \N__35545\
        );

    \I__6422\ : InMux
    port map (
            O => \N__35605\,
            I => \N__35545\
        );

    \I__6421\ : InMux
    port map (
            O => \N__35604\,
            I => \N__35545\
        );

    \I__6420\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35545\
        );

    \I__6419\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35536\
        );

    \I__6418\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35536\
        );

    \I__6417\ : InMux
    port map (
            O => \N__35600\,
            I => \N__35536\
        );

    \I__6416\ : InMux
    port map (
            O => \N__35599\,
            I => \N__35536\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__35590\,
            I => \N__35533\
        );

    \I__6414\ : InMux
    port map (
            O => \N__35589\,
            I => \N__35524\
        );

    \I__6413\ : InMux
    port map (
            O => \N__35588\,
            I => \N__35524\
        );

    \I__6412\ : InMux
    port map (
            O => \N__35587\,
            I => \N__35524\
        );

    \I__6411\ : InMux
    port map (
            O => \N__35586\,
            I => \N__35524\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__35581\,
            I => \N__35519\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__35572\,
            I => \N__35519\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__35563\,
            I => \N__35510\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__35554\,
            I => \N__35510\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__35545\,
            I => \N__35510\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__35536\,
            I => \N__35510\
        );

    \I__6404\ : Span4Mux_h
    port map (
            O => \N__35533\,
            I => \N__35501\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__35524\,
            I => \N__35501\
        );

    \I__6402\ : Span4Mux_v
    port map (
            O => \N__35519\,
            I => \N__35501\
        );

    \I__6401\ : Span4Mux_v
    port map (
            O => \N__35510\,
            I => \N__35501\
        );

    \I__6400\ : Odrv4
    port map (
            O => \N__35501\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6399\ : InMux
    port map (
            O => \N__35498\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__6398\ : InMux
    port map (
            O => \N__35495\,
            I => \N__35491\
        );

    \I__6397\ : InMux
    port map (
            O => \N__35494\,
            I => \N__35488\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__35491\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__35488\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__6394\ : CEMux
    port map (
            O => \N__35483\,
            I => \N__35479\
        );

    \I__6393\ : CEMux
    port map (
            O => \N__35482\,
            I => \N__35476\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__35479\,
            I => \N__35472\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__35476\,
            I => \N__35469\
        );

    \I__6390\ : CEMux
    port map (
            O => \N__35475\,
            I => \N__35466\
        );

    \I__6389\ : Span4Mux_v
    port map (
            O => \N__35472\,
            I => \N__35459\
        );

    \I__6388\ : Span4Mux_v
    port map (
            O => \N__35469\,
            I => \N__35459\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__35466\,
            I => \N__35459\
        );

    \I__6386\ : Span4Mux_v
    port map (
            O => \N__35459\,
            I => \N__35455\
        );

    \I__6385\ : CEMux
    port map (
            O => \N__35458\,
            I => \N__35452\
        );

    \I__6384\ : Span4Mux_v
    port map (
            O => \N__35455\,
            I => \N__35449\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__35452\,
            I => \N__35446\
        );

    \I__6382\ : Odrv4
    port map (
            O => \N__35449\,
            I => \delay_measurement_inst.delay_tr_timer.N_168_i\
        );

    \I__6381\ : Odrv12
    port map (
            O => \N__35446\,
            I => \delay_measurement_inst.delay_tr_timer.N_168_i\
        );

    \I__6380\ : InMux
    port map (
            O => \N__35441\,
            I => \N__35438\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__35438\,
            I => \N__35435\
        );

    \I__6378\ : Span4Mux_v
    port map (
            O => \N__35435\,
            I => \N__35432\
        );

    \I__6377\ : Span4Mux_h
    port map (
            O => \N__35432\,
            I => \N__35429\
        );

    \I__6376\ : Sp12to4
    port map (
            O => \N__35429\,
            I => \N__35426\
        );

    \I__6375\ : Span12Mux_v
    port map (
            O => \N__35426\,
            I => \N__35423\
        );

    \I__6374\ : Odrv12
    port map (
            O => \N__35423\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_0\
        );

    \I__6373\ : CascadeMux
    port map (
            O => \N__35420\,
            I => \N__35417\
        );

    \I__6372\ : InMux
    port map (
            O => \N__35417\,
            I => \N__35414\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__35414\,
            I => \N__35411\
        );

    \I__6370\ : Span4Mux_v
    port map (
            O => \N__35411\,
            I => \N__35408\
        );

    \I__6369\ : Span4Mux_h
    port map (
            O => \N__35408\,
            I => \N__35405\
        );

    \I__6368\ : Sp12to4
    port map (
            O => \N__35405\,
            I => \N__35402\
        );

    \I__6367\ : Odrv12
    port map (
            O => \N__35402\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_15\
        );

    \I__6366\ : InMux
    port map (
            O => \N__35399\,
            I => \N__35396\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__35396\,
            I => \N__35393\
        );

    \I__6364\ : Span4Mux_v
    port map (
            O => \N__35393\,
            I => \N__35390\
        );

    \I__6363\ : Sp12to4
    port map (
            O => \N__35390\,
            I => \N__35387\
        );

    \I__6362\ : Span12Mux_h
    port map (
            O => \N__35387\,
            I => \N__35384\
        );

    \I__6361\ : Odrv12
    port map (
            O => \N__35384\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_16\
        );

    \I__6360\ : CascadeMux
    port map (
            O => \N__35381\,
            I => \N__35378\
        );

    \I__6359\ : InMux
    port map (
            O => \N__35378\,
            I => \N__35375\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__35375\,
            I => \N__35372\
        );

    \I__6357\ : Span12Mux_v
    port map (
            O => \N__35372\,
            I => \N__35369\
        );

    \I__6356\ : Span12Mux_h
    port map (
            O => \N__35369\,
            I => \N__35366\
        );

    \I__6355\ : Odrv12
    port map (
            O => \N__35366\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_1\
        );

    \I__6354\ : InMux
    port map (
            O => \N__35363\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\
        );

    \I__6353\ : InMux
    port map (
            O => \N__35360\,
            I => \N__35357\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__35357\,
            I => \N__35354\
        );

    \I__6351\ : Span4Mux_v
    port map (
            O => \N__35354\,
            I => \N__35351\
        );

    \I__6350\ : Sp12to4
    port map (
            O => \N__35351\,
            I => \N__35348\
        );

    \I__6349\ : Span12Mux_h
    port map (
            O => \N__35348\,
            I => \N__35345\
        );

    \I__6348\ : Odrv12
    port map (
            O => \N__35345\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_17\
        );

    \I__6347\ : CascadeMux
    port map (
            O => \N__35342\,
            I => \N__35339\
        );

    \I__6346\ : InMux
    port map (
            O => \N__35339\,
            I => \N__35336\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__35336\,
            I => \N__35333\
        );

    \I__6344\ : Span12Mux_s10_v
    port map (
            O => \N__35333\,
            I => \N__35330\
        );

    \I__6343\ : Span12Mux_h
    port map (
            O => \N__35330\,
            I => \N__35327\
        );

    \I__6342\ : Odrv12
    port map (
            O => \N__35327\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_2\
        );

    \I__6341\ : InMux
    port map (
            O => \N__35324\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\
        );

    \I__6340\ : InMux
    port map (
            O => \N__35321\,
            I => \N__35318\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__35318\,
            I => \N__35315\
        );

    \I__6338\ : Sp12to4
    port map (
            O => \N__35315\,
            I => \N__35312\
        );

    \I__6337\ : Span12Mux_s9_v
    port map (
            O => \N__35312\,
            I => \N__35309\
        );

    \I__6336\ : Span12Mux_h
    port map (
            O => \N__35309\,
            I => \N__35306\
        );

    \I__6335\ : Odrv12
    port map (
            O => \N__35306\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_3\
        );

    \I__6334\ : CascadeMux
    port map (
            O => \N__35303\,
            I => \N__35300\
        );

    \I__6333\ : InMux
    port map (
            O => \N__35300\,
            I => \N__35297\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__35297\,
            I => \N__35294\
        );

    \I__6331\ : Span4Mux_v
    port map (
            O => \N__35294\,
            I => \N__35291\
        );

    \I__6330\ : Sp12to4
    port map (
            O => \N__35291\,
            I => \N__35288\
        );

    \I__6329\ : Span12Mux_h
    port map (
            O => \N__35288\,
            I => \N__35285\
        );

    \I__6328\ : Odrv12
    port map (
            O => \N__35285\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_18\
        );

    \I__6327\ : InMux
    port map (
            O => \N__35282\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\
        );

    \I__6326\ : InMux
    port map (
            O => \N__35279\,
            I => \N__35276\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__35276\,
            I => \N__35273\
        );

    \I__6324\ : Span12Mux_s8_v
    port map (
            O => \N__35273\,
            I => \N__35270\
        );

    \I__6323\ : Span12Mux_v
    port map (
            O => \N__35270\,
            I => \N__35267\
        );

    \I__6322\ : Odrv12
    port map (
            O => \N__35267\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_4\
        );

    \I__6321\ : InMux
    port map (
            O => \N__35264\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\
        );

    \I__6320\ : CascadeMux
    port map (
            O => \N__35261\,
            I => \N__35258\
        );

    \I__6319\ : InMux
    port map (
            O => \N__35258\,
            I => \N__35253\
        );

    \I__6318\ : InMux
    port map (
            O => \N__35257\,
            I => \N__35250\
        );

    \I__6317\ : InMux
    port map (
            O => \N__35256\,
            I => \N__35247\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__35253\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__35250\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__35247\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__6313\ : InMux
    port map (
            O => \N__35240\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__6312\ : CascadeMux
    port map (
            O => \N__35237\,
            I => \N__35234\
        );

    \I__6311\ : InMux
    port map (
            O => \N__35234\,
            I => \N__35229\
        );

    \I__6310\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35226\
        );

    \I__6309\ : InMux
    port map (
            O => \N__35232\,
            I => \N__35223\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__35229\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__35226\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__35223\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__6305\ : InMux
    port map (
            O => \N__35216\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__6304\ : CascadeMux
    port map (
            O => \N__35213\,
            I => \N__35210\
        );

    \I__6303\ : InMux
    port map (
            O => \N__35210\,
            I => \N__35205\
        );

    \I__6302\ : InMux
    port map (
            O => \N__35209\,
            I => \N__35202\
        );

    \I__6301\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35199\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__35205\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__35202\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__35199\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__6297\ : InMux
    port map (
            O => \N__35192\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__6296\ : CascadeMux
    port map (
            O => \N__35189\,
            I => \N__35186\
        );

    \I__6295\ : InMux
    port map (
            O => \N__35186\,
            I => \N__35181\
        );

    \I__6294\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35178\
        );

    \I__6293\ : InMux
    port map (
            O => \N__35184\,
            I => \N__35175\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__35181\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__35178\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__35175\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__6289\ : InMux
    port map (
            O => \N__35168\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__6288\ : CascadeMux
    port map (
            O => \N__35165\,
            I => \N__35162\
        );

    \I__6287\ : InMux
    port map (
            O => \N__35162\,
            I => \N__35157\
        );

    \I__6286\ : InMux
    port map (
            O => \N__35161\,
            I => \N__35154\
        );

    \I__6285\ : InMux
    port map (
            O => \N__35160\,
            I => \N__35151\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__35157\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__35154\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__35151\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__6281\ : InMux
    port map (
            O => \N__35144\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__6280\ : CascadeMux
    port map (
            O => \N__35141\,
            I => \N__35138\
        );

    \I__6279\ : InMux
    port map (
            O => \N__35138\,
            I => \N__35133\
        );

    \I__6278\ : InMux
    port map (
            O => \N__35137\,
            I => \N__35130\
        );

    \I__6277\ : InMux
    port map (
            O => \N__35136\,
            I => \N__35127\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__35133\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__35130\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__35127\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__6273\ : InMux
    port map (
            O => \N__35120\,
            I => \bfn_12_22_0_\
        );

    \I__6272\ : CascadeMux
    port map (
            O => \N__35117\,
            I => \N__35114\
        );

    \I__6271\ : InMux
    port map (
            O => \N__35114\,
            I => \N__35109\
        );

    \I__6270\ : InMux
    port map (
            O => \N__35113\,
            I => \N__35106\
        );

    \I__6269\ : InMux
    port map (
            O => \N__35112\,
            I => \N__35103\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__35109\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__35106\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__35103\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__6265\ : InMux
    port map (
            O => \N__35096\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__6264\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35088\
        );

    \I__6263\ : InMux
    port map (
            O => \N__35092\,
            I => \N__35083\
        );

    \I__6262\ : InMux
    port map (
            O => \N__35091\,
            I => \N__35083\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__35088\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__35083\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__6259\ : InMux
    port map (
            O => \N__35078\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__6258\ : CascadeMux
    port map (
            O => \N__35075\,
            I => \N__35072\
        );

    \I__6257\ : InMux
    port map (
            O => \N__35072\,
            I => \N__35067\
        );

    \I__6256\ : InMux
    port map (
            O => \N__35071\,
            I => \N__35064\
        );

    \I__6255\ : InMux
    port map (
            O => \N__35070\,
            I => \N__35061\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__35067\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__35064\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__35061\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__6251\ : InMux
    port map (
            O => \N__35054\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__6250\ : CascadeMux
    port map (
            O => \N__35051\,
            I => \N__35048\
        );

    \I__6249\ : InMux
    port map (
            O => \N__35048\,
            I => \N__35043\
        );

    \I__6248\ : InMux
    port map (
            O => \N__35047\,
            I => \N__35040\
        );

    \I__6247\ : InMux
    port map (
            O => \N__35046\,
            I => \N__35037\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__35043\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__35040\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__35037\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__6243\ : InMux
    port map (
            O => \N__35030\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__6242\ : CascadeMux
    port map (
            O => \N__35027\,
            I => \N__35024\
        );

    \I__6241\ : InMux
    port map (
            O => \N__35024\,
            I => \N__35019\
        );

    \I__6240\ : InMux
    port map (
            O => \N__35023\,
            I => \N__35016\
        );

    \I__6239\ : InMux
    port map (
            O => \N__35022\,
            I => \N__35013\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__35019\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__35016\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__35013\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__6235\ : InMux
    port map (
            O => \N__35006\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__6234\ : CascadeMux
    port map (
            O => \N__35003\,
            I => \N__35000\
        );

    \I__6233\ : InMux
    port map (
            O => \N__35000\,
            I => \N__34995\
        );

    \I__6232\ : InMux
    port map (
            O => \N__34999\,
            I => \N__34992\
        );

    \I__6231\ : InMux
    port map (
            O => \N__34998\,
            I => \N__34989\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__34995\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__34992\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__34989\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__6227\ : InMux
    port map (
            O => \N__34982\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__6226\ : CascadeMux
    port map (
            O => \N__34979\,
            I => \N__34976\
        );

    \I__6225\ : InMux
    port map (
            O => \N__34976\,
            I => \N__34971\
        );

    \I__6224\ : InMux
    port map (
            O => \N__34975\,
            I => \N__34968\
        );

    \I__6223\ : InMux
    port map (
            O => \N__34974\,
            I => \N__34965\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__34971\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__34968\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__34965\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__6219\ : InMux
    port map (
            O => \N__34958\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__6218\ : CascadeMux
    port map (
            O => \N__34955\,
            I => \N__34952\
        );

    \I__6217\ : InMux
    port map (
            O => \N__34952\,
            I => \N__34947\
        );

    \I__6216\ : InMux
    port map (
            O => \N__34951\,
            I => \N__34944\
        );

    \I__6215\ : InMux
    port map (
            O => \N__34950\,
            I => \N__34941\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__34947\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__34944\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__34941\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__6211\ : InMux
    port map (
            O => \N__34934\,
            I => \bfn_12_21_0_\
        );

    \I__6210\ : CascadeMux
    port map (
            O => \N__34931\,
            I => \N__34928\
        );

    \I__6209\ : InMux
    port map (
            O => \N__34928\,
            I => \N__34923\
        );

    \I__6208\ : InMux
    port map (
            O => \N__34927\,
            I => \N__34920\
        );

    \I__6207\ : InMux
    port map (
            O => \N__34926\,
            I => \N__34917\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__34923\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__34920\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__34917\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__6203\ : InMux
    port map (
            O => \N__34910\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__6202\ : CascadeMux
    port map (
            O => \N__34907\,
            I => \N__34904\
        );

    \I__6201\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34899\
        );

    \I__6200\ : InMux
    port map (
            O => \N__34903\,
            I => \N__34896\
        );

    \I__6199\ : InMux
    port map (
            O => \N__34902\,
            I => \N__34893\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__34899\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__34896\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__34893\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__6195\ : InMux
    port map (
            O => \N__34886\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__6194\ : InMux
    port map (
            O => \N__34883\,
            I => \N__34878\
        );

    \I__6193\ : InMux
    port map (
            O => \N__34882\,
            I => \N__34873\
        );

    \I__6192\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34873\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__34878\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__34873\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__6189\ : InMux
    port map (
            O => \N__34868\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__6188\ : CascadeMux
    port map (
            O => \N__34865\,
            I => \N__34862\
        );

    \I__6187\ : InMux
    port map (
            O => \N__34862\,
            I => \N__34857\
        );

    \I__6186\ : InMux
    port map (
            O => \N__34861\,
            I => \N__34854\
        );

    \I__6185\ : InMux
    port map (
            O => \N__34860\,
            I => \N__34851\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__34857\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__34854\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__34851\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__6181\ : InMux
    port map (
            O => \N__34844\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__6180\ : CascadeMux
    port map (
            O => \N__34841\,
            I => \N__34836\
        );

    \I__6179\ : CascadeMux
    port map (
            O => \N__34840\,
            I => \N__34833\
        );

    \I__6178\ : InMux
    port map (
            O => \N__34839\,
            I => \N__34830\
        );

    \I__6177\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34825\
        );

    \I__6176\ : InMux
    port map (
            O => \N__34833\,
            I => \N__34825\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__34830\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__34825\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__6173\ : InMux
    port map (
            O => \N__34820\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__34817\,
            I => \N__34814\
        );

    \I__6171\ : InMux
    port map (
            O => \N__34814\,
            I => \N__34809\
        );

    \I__6170\ : InMux
    port map (
            O => \N__34813\,
            I => \N__34806\
        );

    \I__6169\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34803\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__34809\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__34806\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__34803\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__6165\ : InMux
    port map (
            O => \N__34796\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__6164\ : CascadeMux
    port map (
            O => \N__34793\,
            I => \N__34790\
        );

    \I__6163\ : InMux
    port map (
            O => \N__34790\,
            I => \N__34785\
        );

    \I__6162\ : InMux
    port map (
            O => \N__34789\,
            I => \N__34782\
        );

    \I__6161\ : InMux
    port map (
            O => \N__34788\,
            I => \N__34779\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__34785\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__34782\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__34779\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__6157\ : InMux
    port map (
            O => \N__34772\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__6156\ : CascadeMux
    port map (
            O => \N__34769\,
            I => \N__34766\
        );

    \I__6155\ : InMux
    port map (
            O => \N__34766\,
            I => \N__34761\
        );

    \I__6154\ : InMux
    port map (
            O => \N__34765\,
            I => \N__34758\
        );

    \I__6153\ : InMux
    port map (
            O => \N__34764\,
            I => \N__34755\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__34761\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__34758\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__34755\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__6149\ : InMux
    port map (
            O => \N__34748\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__6148\ : CascadeMux
    port map (
            O => \N__34745\,
            I => \N__34742\
        );

    \I__6147\ : InMux
    port map (
            O => \N__34742\,
            I => \N__34737\
        );

    \I__6146\ : InMux
    port map (
            O => \N__34741\,
            I => \N__34734\
        );

    \I__6145\ : InMux
    port map (
            O => \N__34740\,
            I => \N__34731\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__34737\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__34734\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__34731\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__6141\ : InMux
    port map (
            O => \N__34724\,
            I => \bfn_12_20_0_\
        );

    \I__6140\ : CascadeMux
    port map (
            O => \N__34721\,
            I => \N__34718\
        );

    \I__6139\ : InMux
    port map (
            O => \N__34718\,
            I => \N__34713\
        );

    \I__6138\ : InMux
    port map (
            O => \N__34717\,
            I => \N__34710\
        );

    \I__6137\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34707\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__34713\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__34710\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__34707\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__6133\ : InMux
    port map (
            O => \N__34700\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__6132\ : CascadeMux
    port map (
            O => \N__34697\,
            I => \N__34694\
        );

    \I__6131\ : InMux
    port map (
            O => \N__34694\,
            I => \N__34689\
        );

    \I__6130\ : InMux
    port map (
            O => \N__34693\,
            I => \N__34686\
        );

    \I__6129\ : InMux
    port map (
            O => \N__34692\,
            I => \N__34683\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__34689\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__34686\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__34683\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__6125\ : InMux
    port map (
            O => \N__34676\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__6124\ : InMux
    port map (
            O => \N__34673\,
            I => \N__34670\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__34670\,
            I => \N__34666\
        );

    \I__6122\ : InMux
    port map (
            O => \N__34669\,
            I => \N__34663\
        );

    \I__6121\ : Odrv12
    port map (
            O => \N__34666\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_17
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__34663\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_17
        );

    \I__6119\ : InMux
    port map (
            O => \N__34658\,
            I => \N__34652\
        );

    \I__6118\ : InMux
    port map (
            O => \N__34657\,
            I => \N__34652\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__34652\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_17\
        );

    \I__6116\ : InMux
    port map (
            O => \N__34649\,
            I => \N__34646\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__34646\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt18\
        );

    \I__6114\ : InMux
    port map (
            O => \N__34643\,
            I => \N__34639\
        );

    \I__6113\ : InMux
    port map (
            O => \N__34642\,
            I => \N__34636\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__34639\,
            I => \N__34633\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__34636\,
            I => \N__34630\
        );

    \I__6110\ : Odrv12
    port map (
            O => \N__34633\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_18
        );

    \I__6109\ : Odrv4
    port map (
            O => \N__34630\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_18
        );

    \I__6108\ : InMux
    port map (
            O => \N__34625\,
            I => \N__34619\
        );

    \I__6107\ : InMux
    port map (
            O => \N__34624\,
            I => \N__34619\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__34619\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_18\
        );

    \I__6105\ : InMux
    port map (
            O => \N__34616\,
            I => \N__34610\
        );

    \I__6104\ : InMux
    port map (
            O => \N__34615\,
            I => \N__34610\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__34610\,
            I => \N__34607\
        );

    \I__6102\ : Odrv4
    port map (
            O => \N__34607\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_19\
        );

    \I__6101\ : CascadeMux
    port map (
            O => \N__34604\,
            I => \N__34600\
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__34603\,
            I => \N__34597\
        );

    \I__6099\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34592\
        );

    \I__6098\ : InMux
    port map (
            O => \N__34597\,
            I => \N__34592\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__34592\,
            I => \N__34588\
        );

    \I__6096\ : InMux
    port map (
            O => \N__34591\,
            I => \N__34585\
        );

    \I__6095\ : Span4Mux_h
    port map (
            O => \N__34588\,
            I => \N__34582\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__34585\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_19\
        );

    \I__6093\ : Odrv4
    port map (
            O => \N__34582\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_19\
        );

    \I__6092\ : InMux
    port map (
            O => \N__34577\,
            I => \N__34571\
        );

    \I__6091\ : InMux
    port map (
            O => \N__34576\,
            I => \N__34571\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__34571\,
            I => \N__34567\
        );

    \I__6089\ : InMux
    port map (
            O => \N__34570\,
            I => \N__34564\
        );

    \I__6088\ : Span4Mux_h
    port map (
            O => \N__34567\,
            I => \N__34561\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__34564\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_18\
        );

    \I__6086\ : Odrv4
    port map (
            O => \N__34561\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_18\
        );

    \I__6085\ : CascadeMux
    port map (
            O => \N__34556\,
            I => \N__34553\
        );

    \I__6084\ : InMux
    port map (
            O => \N__34553\,
            I => \N__34550\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__34550\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18\
        );

    \I__6082\ : CascadeMux
    port map (
            O => \N__34547\,
            I => \N__34540\
        );

    \I__6081\ : InMux
    port map (
            O => \N__34546\,
            I => \N__34537\
        );

    \I__6080\ : InMux
    port map (
            O => \N__34545\,
            I => \N__34534\
        );

    \I__6079\ : InMux
    port map (
            O => \N__34544\,
            I => \N__34531\
        );

    \I__6078\ : InMux
    port map (
            O => \N__34543\,
            I => \N__34528\
        );

    \I__6077\ : InMux
    port map (
            O => \N__34540\,
            I => \N__34524\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__34537\,
            I => \N__34517\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__34534\,
            I => \N__34517\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__34531\,
            I => \N__34517\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__34528\,
            I => \N__34514\
        );

    \I__6072\ : InMux
    port map (
            O => \N__34527\,
            I => \N__34511\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__34524\,
            I => \N__34506\
        );

    \I__6070\ : Span4Mux_v
    port map (
            O => \N__34517\,
            I => \N__34506\
        );

    \I__6069\ : Span4Mux_v
    port map (
            O => \N__34514\,
            I => \N__34503\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__34511\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__6067\ : Odrv4
    port map (
            O => \N__34506\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__6066\ : Odrv4
    port map (
            O => \N__34503\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__6065\ : InMux
    port map (
            O => \N__34496\,
            I => \N__34472\
        );

    \I__6064\ : InMux
    port map (
            O => \N__34495\,
            I => \N__34472\
        );

    \I__6063\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34472\
        );

    \I__6062\ : InMux
    port map (
            O => \N__34493\,
            I => \N__34472\
        );

    \I__6061\ : InMux
    port map (
            O => \N__34492\,
            I => \N__34463\
        );

    \I__6060\ : InMux
    port map (
            O => \N__34491\,
            I => \N__34463\
        );

    \I__6059\ : InMux
    port map (
            O => \N__34490\,
            I => \N__34463\
        );

    \I__6058\ : InMux
    port map (
            O => \N__34489\,
            I => \N__34463\
        );

    \I__6057\ : InMux
    port map (
            O => \N__34488\,
            I => \N__34446\
        );

    \I__6056\ : InMux
    port map (
            O => \N__34487\,
            I => \N__34446\
        );

    \I__6055\ : InMux
    port map (
            O => \N__34486\,
            I => \N__34446\
        );

    \I__6054\ : InMux
    port map (
            O => \N__34485\,
            I => \N__34446\
        );

    \I__6053\ : InMux
    port map (
            O => \N__34484\,
            I => \N__34437\
        );

    \I__6052\ : InMux
    port map (
            O => \N__34483\,
            I => \N__34437\
        );

    \I__6051\ : InMux
    port map (
            O => \N__34482\,
            I => \N__34437\
        );

    \I__6050\ : InMux
    port map (
            O => \N__34481\,
            I => \N__34437\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__34472\,
            I => \N__34428\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__34463\,
            I => \N__34428\
        );

    \I__6047\ : InMux
    port map (
            O => \N__34462\,
            I => \N__34421\
        );

    \I__6046\ : InMux
    port map (
            O => \N__34461\,
            I => \N__34421\
        );

    \I__6045\ : InMux
    port map (
            O => \N__34460\,
            I => \N__34421\
        );

    \I__6044\ : InMux
    port map (
            O => \N__34459\,
            I => \N__34410\
        );

    \I__6043\ : InMux
    port map (
            O => \N__34458\,
            I => \N__34410\
        );

    \I__6042\ : InMux
    port map (
            O => \N__34457\,
            I => \N__34410\
        );

    \I__6041\ : InMux
    port map (
            O => \N__34456\,
            I => \N__34410\
        );

    \I__6040\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34410\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__34446\,
            I => \N__34401\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__34437\,
            I => \N__34401\
        );

    \I__6037\ : InMux
    port map (
            O => \N__34436\,
            I => \N__34392\
        );

    \I__6036\ : InMux
    port map (
            O => \N__34435\,
            I => \N__34392\
        );

    \I__6035\ : InMux
    port map (
            O => \N__34434\,
            I => \N__34392\
        );

    \I__6034\ : InMux
    port map (
            O => \N__34433\,
            I => \N__34392\
        );

    \I__6033\ : Span4Mux_v
    port map (
            O => \N__34428\,
            I => \N__34387\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__34421\,
            I => \N__34387\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__34410\,
            I => \N__34384\
        );

    \I__6030\ : InMux
    port map (
            O => \N__34409\,
            I => \N__34375\
        );

    \I__6029\ : InMux
    port map (
            O => \N__34408\,
            I => \N__34375\
        );

    \I__6028\ : InMux
    port map (
            O => \N__34407\,
            I => \N__34375\
        );

    \I__6027\ : InMux
    port map (
            O => \N__34406\,
            I => \N__34375\
        );

    \I__6026\ : Span4Mux_h
    port map (
            O => \N__34401\,
            I => \N__34366\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__34392\,
            I => \N__34366\
        );

    \I__6024\ : Span4Mux_v
    port map (
            O => \N__34387\,
            I => \N__34366\
        );

    \I__6023\ : Span4Mux_v
    port map (
            O => \N__34384\,
            I => \N__34366\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__34375\,
            I => \phase_controller_inst1.stoper_hc.start_latched_i_0\
        );

    \I__6021\ : Odrv4
    port map (
            O => \N__34366\,
            I => \phase_controller_inst1.stoper_hc.start_latched_i_0\
        );

    \I__6020\ : InMux
    port map (
            O => \N__34361\,
            I => \N__34355\
        );

    \I__6019\ : InMux
    port map (
            O => \N__34360\,
            I => \N__34348\
        );

    \I__6018\ : InMux
    port map (
            O => \N__34359\,
            I => \N__34348\
        );

    \I__6017\ : InMux
    port map (
            O => \N__34358\,
            I => \N__34348\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__34355\,
            I => \N__34345\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__34348\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6014\ : Odrv12
    port map (
            O => \N__34345\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6013\ : InMux
    port map (
            O => \N__34340\,
            I => \N__34337\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__34337\,
            I => \N__34334\
        );

    \I__6011\ : Span4Mux_h
    port map (
            O => \N__34334\,
            I => \N__34330\
        );

    \I__6010\ : CascadeMux
    port map (
            O => \N__34333\,
            I => \N__34327\
        );

    \I__6009\ : Span4Mux_v
    port map (
            O => \N__34330\,
            I => \N__34323\
        );

    \I__6008\ : InMux
    port map (
            O => \N__34327\,
            I => \N__34320\
        );

    \I__6007\ : InMux
    port map (
            O => \N__34326\,
            I => \N__34317\
        );

    \I__6006\ : Odrv4
    port map (
            O => \N__34323\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__34320\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__34317\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__6003\ : InMux
    port map (
            O => \N__34310\,
            I => \bfn_12_19_0_\
        );

    \I__6002\ : InMux
    port map (
            O => \N__34307\,
            I => \N__34304\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__34304\,
            I => \N__34301\
        );

    \I__6000\ : Span4Mux_v
    port map (
            O => \N__34301\,
            I => \N__34298\
        );

    \I__5999\ : Span4Mux_v
    port map (
            O => \N__34298\,
            I => \N__34294\
        );

    \I__5998\ : CascadeMux
    port map (
            O => \N__34297\,
            I => \N__34291\
        );

    \I__5997\ : Span4Mux_h
    port map (
            O => \N__34294\,
            I => \N__34287\
        );

    \I__5996\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34284\
        );

    \I__5995\ : InMux
    port map (
            O => \N__34290\,
            I => \N__34281\
        );

    \I__5994\ : Odrv4
    port map (
            O => \N__34287\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__34284\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__34281\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__5991\ : InMux
    port map (
            O => \N__34274\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__5990\ : CEMux
    port map (
            O => \N__34271\,
            I => \N__34266\
        );

    \I__5989\ : CEMux
    port map (
            O => \N__34270\,
            I => \N__34263\
        );

    \I__5988\ : CEMux
    port map (
            O => \N__34269\,
            I => \N__34260\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__34266\,
            I => \N__34256\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__34263\,
            I => \N__34251\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__34260\,
            I => \N__34251\
        );

    \I__5984\ : CEMux
    port map (
            O => \N__34259\,
            I => \N__34248\
        );

    \I__5983\ : Span4Mux_v
    port map (
            O => \N__34256\,
            I => \N__34241\
        );

    \I__5982\ : Span4Mux_v
    port map (
            O => \N__34251\,
            I => \N__34241\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__34248\,
            I => \N__34238\
        );

    \I__5980\ : CEMux
    port map (
            O => \N__34247\,
            I => \N__34235\
        );

    \I__5979\ : CEMux
    port map (
            O => \N__34246\,
            I => \N__34232\
        );

    \I__5978\ : Span4Mux_v
    port map (
            O => \N__34241\,
            I => \N__34227\
        );

    \I__5977\ : Span4Mux_v
    port map (
            O => \N__34238\,
            I => \N__34227\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__34235\,
            I => \N__34224\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__34232\,
            I => \N__34221\
        );

    \I__5974\ : Span4Mux_v
    port map (
            O => \N__34227\,
            I => \N__34218\
        );

    \I__5973\ : Span4Mux_v
    port map (
            O => \N__34224\,
            I => \N__34215\
        );

    \I__5972\ : Span4Mux_h
    port map (
            O => \N__34221\,
            I => \N__34212\
        );

    \I__5971\ : Odrv4
    port map (
            O => \N__34218\,
            I => \delay_measurement_inst.delay_tr_timer.N_167_i\
        );

    \I__5970\ : Odrv4
    port map (
            O => \N__34215\,
            I => \delay_measurement_inst.delay_tr_timer.N_167_i\
        );

    \I__5969\ : Odrv4
    port map (
            O => \N__34212\,
            I => \delay_measurement_inst.delay_tr_timer.N_167_i\
        );

    \I__5968\ : InMux
    port map (
            O => \N__34205\,
            I => \N__34202\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__34202\,
            I => \N__34199\
        );

    \I__5966\ : Span4Mux_h
    port map (
            O => \N__34199\,
            I => \N__34194\
        );

    \I__5965\ : InMux
    port map (
            O => \N__34198\,
            I => \N__34191\
        );

    \I__5964\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34188\
        );

    \I__5963\ : Odrv4
    port map (
            O => \N__34194\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__34191\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__34188\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__5960\ : CascadeMux
    port map (
            O => \N__34181\,
            I => \phase_controller_inst1.stoper_hc.un4_start_0_cascade_\
        );

    \I__5959\ : InMux
    port map (
            O => \N__34178\,
            I => \N__34175\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__34175\,
            I => \N__34171\
        );

    \I__5957\ : InMux
    port map (
            O => \N__34174\,
            I => \N__34168\
        );

    \I__5956\ : Span4Mux_h
    port map (
            O => \N__34171\,
            I => \N__34162\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__34168\,
            I => \N__34162\
        );

    \I__5954\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34159\
        );

    \I__5953\ : Odrv4
    port map (
            O => \N__34162\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__34159\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO\
        );

    \I__5951\ : CascadeMux
    port map (
            O => \N__34154\,
            I => \N__34150\
        );

    \I__5950\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34145\
        );

    \I__5949\ : InMux
    port map (
            O => \N__34150\,
            I => \N__34145\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__34145\,
            I => \N__34140\
        );

    \I__5947\ : InMux
    port map (
            O => \N__34144\,
            I => \N__34137\
        );

    \I__5946\ : InMux
    port map (
            O => \N__34143\,
            I => \N__34134\
        );

    \I__5945\ : Span4Mux_v
    port map (
            O => \N__34140\,
            I => \N__34129\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__34137\,
            I => \N__34129\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__34134\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5942\ : Odrv4
    port map (
            O => \N__34129\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5941\ : InMux
    port map (
            O => \N__34124\,
            I => \N__34120\
        );

    \I__5940\ : InMux
    port map (
            O => \N__34123\,
            I => \N__34117\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__34120\,
            I => \N__34113\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__34117\,
            I => \N__34110\
        );

    \I__5937\ : InMux
    port map (
            O => \N__34116\,
            I => \N__34107\
        );

    \I__5936\ : Span4Mux_v
    port map (
            O => \N__34113\,
            I => \N__34102\
        );

    \I__5935\ : Span4Mux_h
    port map (
            O => \N__34110\,
            I => \N__34102\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__34107\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_31\
        );

    \I__5933\ : Odrv4
    port map (
            O => \N__34102\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_31\
        );

    \I__5932\ : InMux
    port map (
            O => \N__34097\,
            I => \N__34094\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__34094\,
            I => \N__34090\
        );

    \I__5930\ : InMux
    port map (
            O => \N__34093\,
            I => \N__34087\
        );

    \I__5929\ : Span4Mux_v
    port map (
            O => \N__34090\,
            I => \N__34081\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__34087\,
            I => \N__34081\
        );

    \I__5927\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34078\
        );

    \I__5926\ : Span4Mux_h
    port map (
            O => \N__34081\,
            I => \N__34075\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__34078\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_30\
        );

    \I__5924\ : Odrv4
    port map (
            O => \N__34075\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_30\
        );

    \I__5923\ : InMux
    port map (
            O => \N__34070\,
            I => \N__34067\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__34067\,
            I => \N__34064\
        );

    \I__5921\ : Span4Mux_v
    port map (
            O => \N__34064\,
            I => \N__34058\
        );

    \I__5920\ : InMux
    port map (
            O => \N__34063\,
            I => \N__34051\
        );

    \I__5919\ : InMux
    port map (
            O => \N__34062\,
            I => \N__34051\
        );

    \I__5918\ : InMux
    port map (
            O => \N__34061\,
            I => \N__34051\
        );

    \I__5917\ : Span4Mux_h
    port map (
            O => \N__34058\,
            I => \N__34046\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__34051\,
            I => \N__34046\
        );

    \I__5915\ : Odrv4
    port map (
            O => \N__34046\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28\
        );

    \I__5914\ : InMux
    port map (
            O => \N__34043\,
            I => \N__34040\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__34040\,
            I => \N__34037\
        );

    \I__5912\ : Span4Mux_h
    port map (
            O => \N__34037\,
            I => \N__34034\
        );

    \I__5911\ : Odrv4
    port map (
            O => \N__34034\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30\
        );

    \I__5910\ : InMux
    port map (
            O => \N__34031\,
            I => \N__34027\
        );

    \I__5909\ : InMux
    port map (
            O => \N__34030\,
            I => \N__34024\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__34027\,
            I => \N__34018\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__34024\,
            I => \N__34014\
        );

    \I__5906\ : InMux
    port map (
            O => \N__34023\,
            I => \N__34007\
        );

    \I__5905\ : InMux
    port map (
            O => \N__34022\,
            I => \N__34007\
        );

    \I__5904\ : InMux
    port map (
            O => \N__34021\,
            I => \N__34007\
        );

    \I__5903\ : Span4Mux_v
    port map (
            O => \N__34018\,
            I => \N__34004\
        );

    \I__5902\ : InMux
    port map (
            O => \N__34017\,
            I => \N__34001\
        );

    \I__5901\ : Span4Mux_h
    port map (
            O => \N__34014\,
            I => \N__33998\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__34007\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5899\ : Odrv4
    port map (
            O => \N__34004\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__34001\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__33998\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5896\ : InMux
    port map (
            O => \N__33989\,
            I => \N__33986\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__33986\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt16\
        );

    \I__5894\ : InMux
    port map (
            O => \N__33983\,
            I => \N__33979\
        );

    \I__5893\ : InMux
    port map (
            O => \N__33982\,
            I => \N__33976\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__33979\,
            I => \N__33973\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__33976\,
            I => \N__33970\
        );

    \I__5890\ : Odrv12
    port map (
            O => \N__33973\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_16
        );

    \I__5889\ : Odrv4
    port map (
            O => \N__33970\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_16
        );

    \I__5888\ : InMux
    port map (
            O => \N__33965\,
            I => \N__33959\
        );

    \I__5887\ : InMux
    port map (
            O => \N__33964\,
            I => \N__33959\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__33959\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_16\
        );

    \I__5885\ : InMux
    port map (
            O => \N__33956\,
            I => \N__33950\
        );

    \I__5884\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33950\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__33950\,
            I => \N__33946\
        );

    \I__5882\ : InMux
    port map (
            O => \N__33949\,
            I => \N__33943\
        );

    \I__5881\ : Span4Mux_h
    port map (
            O => \N__33946\,
            I => \N__33940\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__33943\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_17\
        );

    \I__5879\ : Odrv4
    port map (
            O => \N__33940\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_17\
        );

    \I__5878\ : CascadeMux
    port map (
            O => \N__33935\,
            I => \N__33931\
        );

    \I__5877\ : CascadeMux
    port map (
            O => \N__33934\,
            I => \N__33928\
        );

    \I__5876\ : InMux
    port map (
            O => \N__33931\,
            I => \N__33923\
        );

    \I__5875\ : InMux
    port map (
            O => \N__33928\,
            I => \N__33923\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__33923\,
            I => \N__33919\
        );

    \I__5873\ : InMux
    port map (
            O => \N__33922\,
            I => \N__33916\
        );

    \I__5872\ : Span4Mux_h
    port map (
            O => \N__33919\,
            I => \N__33913\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__33916\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_16\
        );

    \I__5870\ : Odrv4
    port map (
            O => \N__33913\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_16\
        );

    \I__5869\ : CascadeMux
    port map (
            O => \N__33908\,
            I => \N__33905\
        );

    \I__5868\ : InMux
    port map (
            O => \N__33905\,
            I => \N__33902\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__33902\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16\
        );

    \I__5866\ : InMux
    port map (
            O => \N__33899\,
            I => \N__33896\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__33896\,
            I => \N__33892\
        );

    \I__5864\ : InMux
    port map (
            O => \N__33895\,
            I => \N__33889\
        );

    \I__5863\ : Span4Mux_v
    port map (
            O => \N__33892\,
            I => \N__33884\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__33889\,
            I => \N__33884\
        );

    \I__5861\ : Odrv4
    port map (
            O => \N__33884\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_2
        );

    \I__5860\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33878\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__33878\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_2\
        );

    \I__5858\ : InMux
    port map (
            O => \N__33875\,
            I => \N__33871\
        );

    \I__5857\ : InMux
    port map (
            O => \N__33874\,
            I => \N__33868\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__33871\,
            I => \N__33865\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__33868\,
            I => \N__33862\
        );

    \I__5854\ : Odrv12
    port map (
            O => \N__33865\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_6
        );

    \I__5853\ : Odrv4
    port map (
            O => \N__33862\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_6
        );

    \I__5852\ : CascadeMux
    port map (
            O => \N__33857\,
            I => \N__33854\
        );

    \I__5851\ : InMux
    port map (
            O => \N__33854\,
            I => \N__33851\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__33851\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_6\
        );

    \I__5849\ : InMux
    port map (
            O => \N__33848\,
            I => \N__33845\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__33845\,
            I => \N__33841\
        );

    \I__5847\ : InMux
    port map (
            O => \N__33844\,
            I => \N__33838\
        );

    \I__5846\ : Odrv4
    port map (
            O => \N__33841\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_19
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__33838\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_19
        );

    \I__5844\ : InMux
    port map (
            O => \N__33833\,
            I => \N__33830\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__33830\,
            I => \N__33826\
        );

    \I__5842\ : InMux
    port map (
            O => \N__33829\,
            I => \N__33823\
        );

    \I__5841\ : Span4Mux_v
    port map (
            O => \N__33826\,
            I => \N__33818\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__33823\,
            I => \N__33818\
        );

    \I__5839\ : Odrv4
    port map (
            O => \N__33818\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_3
        );

    \I__5838\ : InMux
    port map (
            O => \N__33815\,
            I => \N__33812\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__33812\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_3\
        );

    \I__5836\ : InMux
    port map (
            O => \N__33809\,
            I => \N__33805\
        );

    \I__5835\ : InMux
    port map (
            O => \N__33808\,
            I => \N__33802\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__33805\,
            I => \N__33799\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__33802\,
            I => \N__33796\
        );

    \I__5832\ : Odrv12
    port map (
            O => \N__33799\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_7
        );

    \I__5831\ : Odrv4
    port map (
            O => \N__33796\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_7
        );

    \I__5830\ : CascadeMux
    port map (
            O => \N__33791\,
            I => \N__33788\
        );

    \I__5829\ : InMux
    port map (
            O => \N__33788\,
            I => \N__33785\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__33785\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_7\
        );

    \I__5827\ : InMux
    port map (
            O => \N__33782\,
            I => \N__33778\
        );

    \I__5826\ : InMux
    port map (
            O => \N__33781\,
            I => \N__33775\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__33778\,
            I => \N__33772\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__33775\,
            I => \N__33769\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__33772\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_10
        );

    \I__5822\ : Odrv4
    port map (
            O => \N__33769\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_10
        );

    \I__5821\ : InMux
    port map (
            O => \N__33764\,
            I => \N__33761\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__33761\,
            I => \N__33758\
        );

    \I__5819\ : Odrv4
    port map (
            O => \N__33758\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_10\
        );

    \I__5818\ : InMux
    port map (
            O => \N__33755\,
            I => \N__33751\
        );

    \I__5817\ : InMux
    port map (
            O => \N__33754\,
            I => \N__33748\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__33751\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_25
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__33748\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_25
        );

    \I__5814\ : InMux
    port map (
            O => \N__33743\,
            I => \N__33737\
        );

    \I__5813\ : InMux
    port map (
            O => \N__33742\,
            I => \N__33737\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__33737\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25\
        );

    \I__5811\ : InMux
    port map (
            O => \N__33734\,
            I => \N__33730\
        );

    \I__5810\ : InMux
    port map (
            O => \N__33733\,
            I => \N__33727\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__33730\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_22
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__33727\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_22
        );

    \I__5807\ : InMux
    port map (
            O => \N__33722\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21\
        );

    \I__5806\ : InMux
    port map (
            O => \N__33719\,
            I => \N__33715\
        );

    \I__5805\ : InMux
    port map (
            O => \N__33718\,
            I => \N__33712\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__33715\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_23
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__33712\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_23
        );

    \I__5802\ : InMux
    port map (
            O => \N__33707\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22\
        );

    \I__5801\ : InMux
    port map (
            O => \N__33704\,
            I => \N__33700\
        );

    \I__5800\ : InMux
    port map (
            O => \N__33703\,
            I => \N__33697\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__33700\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_24
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__33697\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_24
        );

    \I__5797\ : InMux
    port map (
            O => \N__33692\,
            I => \bfn_12_10_0_\
        );

    \I__5796\ : InMux
    port map (
            O => \N__33689\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24\
        );

    \I__5795\ : InMux
    port map (
            O => \N__33686\,
            I => \N__33682\
        );

    \I__5794\ : InMux
    port map (
            O => \N__33685\,
            I => \N__33679\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__33682\,
            I => \N__33676\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__33679\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_26
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__33676\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_26
        );

    \I__5790\ : InMux
    port map (
            O => \N__33671\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25\
        );

    \I__5789\ : InMux
    port map (
            O => \N__33668\,
            I => \N__33664\
        );

    \I__5788\ : InMux
    port map (
            O => \N__33667\,
            I => \N__33661\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__33664\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_27
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__33661\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_27
        );

    \I__5785\ : InMux
    port map (
            O => \N__33656\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26\
        );

    \I__5784\ : InMux
    port map (
            O => \N__33653\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27\
        );

    \I__5783\ : InMux
    port map (
            O => \N__33650\,
            I => \N__33646\
        );

    \I__5782\ : InMux
    port map (
            O => \N__33649\,
            I => \N__33643\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__33646\,
            I => \N__33640\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__33643\,
            I => \N__33637\
        );

    \I__5779\ : Odrv12
    port map (
            O => \N__33640\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_4
        );

    \I__5778\ : Odrv4
    port map (
            O => \N__33637\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_4
        );

    \I__5777\ : InMux
    port map (
            O => \N__33632\,
            I => \N__33629\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__33629\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_4\
        );

    \I__5775\ : InMux
    port map (
            O => \N__33626\,
            I => \N__33623\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__33623\,
            I => \N__33619\
        );

    \I__5773\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33616\
        );

    \I__5772\ : Odrv4
    port map (
            O => \N__33619\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_13
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__33616\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_13
        );

    \I__5770\ : InMux
    port map (
            O => \N__33611\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12\
        );

    \I__5769\ : InMux
    port map (
            O => \N__33608\,
            I => \N__33605\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__33605\,
            I => \N__33601\
        );

    \I__5767\ : InMux
    port map (
            O => \N__33604\,
            I => \N__33598\
        );

    \I__5766\ : Odrv4
    port map (
            O => \N__33601\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_14
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__33598\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_14
        );

    \I__5764\ : InMux
    port map (
            O => \N__33593\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13\
        );

    \I__5763\ : InMux
    port map (
            O => \N__33590\,
            I => \N__33587\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__33587\,
            I => \N__33583\
        );

    \I__5761\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33580\
        );

    \I__5760\ : Odrv4
    port map (
            O => \N__33583\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_15
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__33580\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_15
        );

    \I__5758\ : InMux
    port map (
            O => \N__33575\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14\
        );

    \I__5757\ : InMux
    port map (
            O => \N__33572\,
            I => \bfn_12_9_0_\
        );

    \I__5756\ : InMux
    port map (
            O => \N__33569\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16\
        );

    \I__5755\ : InMux
    port map (
            O => \N__33566\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17\
        );

    \I__5754\ : InMux
    port map (
            O => \N__33563\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18\
        );

    \I__5753\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33556\
        );

    \I__5752\ : InMux
    port map (
            O => \N__33559\,
            I => \N__33553\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__33556\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_20
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__33553\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_20
        );

    \I__5749\ : InMux
    port map (
            O => \N__33548\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19\
        );

    \I__5748\ : InMux
    port map (
            O => \N__33545\,
            I => \N__33542\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__33542\,
            I => \N__33538\
        );

    \I__5746\ : InMux
    port map (
            O => \N__33541\,
            I => \N__33535\
        );

    \I__5745\ : Odrv4
    port map (
            O => \N__33538\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_21
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__33535\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_21
        );

    \I__5743\ : InMux
    port map (
            O => \N__33530\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20\
        );

    \I__5742\ : InMux
    port map (
            O => \N__33527\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3\
        );

    \I__5741\ : InMux
    port map (
            O => \N__33524\,
            I => \N__33521\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__33521\,
            I => \N__33517\
        );

    \I__5739\ : InMux
    port map (
            O => \N__33520\,
            I => \N__33514\
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__33517\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_5
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__33514\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_5
        );

    \I__5736\ : InMux
    port map (
            O => \N__33509\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4\
        );

    \I__5735\ : InMux
    port map (
            O => \N__33506\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5\
        );

    \I__5734\ : InMux
    port map (
            O => \N__33503\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6\
        );

    \I__5733\ : InMux
    port map (
            O => \N__33500\,
            I => \N__33497\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__33497\,
            I => \N__33493\
        );

    \I__5731\ : InMux
    port map (
            O => \N__33496\,
            I => \N__33490\
        );

    \I__5730\ : Odrv4
    port map (
            O => \N__33493\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_8
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__33490\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_8
        );

    \I__5728\ : InMux
    port map (
            O => \N__33485\,
            I => \bfn_12_8_0_\
        );

    \I__5727\ : InMux
    port map (
            O => \N__33482\,
            I => \N__33479\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__33479\,
            I => \N__33475\
        );

    \I__5725\ : InMux
    port map (
            O => \N__33478\,
            I => \N__33472\
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__33475\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_9
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__33472\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_9
        );

    \I__5722\ : InMux
    port map (
            O => \N__33467\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8\
        );

    \I__5721\ : InMux
    port map (
            O => \N__33464\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9\
        );

    \I__5720\ : InMux
    port map (
            O => \N__33461\,
            I => \N__33457\
        );

    \I__5719\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33454\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__33457\,
            I => \N__33451\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__33454\,
            I => \N__33448\
        );

    \I__5716\ : Odrv4
    port map (
            O => \N__33451\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_11
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__33448\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_11
        );

    \I__5714\ : InMux
    port map (
            O => \N__33443\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10\
        );

    \I__5713\ : InMux
    port map (
            O => \N__33440\,
            I => \N__33437\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__33437\,
            I => \N__33433\
        );

    \I__5711\ : InMux
    port map (
            O => \N__33436\,
            I => \N__33430\
        );

    \I__5710\ : Odrv4
    port map (
            O => \N__33433\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_12
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__33430\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_12
        );

    \I__5708\ : InMux
    port map (
            O => \N__33425\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11\
        );

    \I__5707\ : InMux
    port map (
            O => \N__33422\,
            I => \N__33419\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__33419\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_14\
        );

    \I__5705\ : InMux
    port map (
            O => \N__33416\,
            I => \N__33413\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__33413\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_13\
        );

    \I__5703\ : InMux
    port map (
            O => \N__33410\,
            I => \N__33407\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__33407\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_8\
        );

    \I__5701\ : CascadeMux
    port map (
            O => \N__33404\,
            I => \N__33401\
        );

    \I__5700\ : InMux
    port map (
            O => \N__33401\,
            I => \N__33398\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__33398\,
            I => \N__33395\
        );

    \I__5698\ : Span4Mux_h
    port map (
            O => \N__33395\,
            I => \N__33392\
        );

    \I__5697\ : Odrv4
    port map (
            O => \N__33392\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_0\
        );

    \I__5696\ : CascadeMux
    port map (
            O => \N__33389\,
            I => \N__33386\
        );

    \I__5695\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33383\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__33383\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_15\
        );

    \I__5693\ : CEMux
    port map (
            O => \N__33380\,
            I => \N__33377\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__33377\,
            I => \N__33371\
        );

    \I__5691\ : CEMux
    port map (
            O => \N__33376\,
            I => \N__33368\
        );

    \I__5690\ : CEMux
    port map (
            O => \N__33375\,
            I => \N__33364\
        );

    \I__5689\ : CEMux
    port map (
            O => \N__33374\,
            I => \N__33361\
        );

    \I__5688\ : Span4Mux_h
    port map (
            O => \N__33371\,
            I => \N__33356\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__33368\,
            I => \N__33356\
        );

    \I__5686\ : CEMux
    port map (
            O => \N__33367\,
            I => \N__33353\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__33364\,
            I => \N__33349\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__33361\,
            I => \N__33346\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__33356\,
            I => \N__33341\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__33353\,
            I => \N__33341\
        );

    \I__5681\ : CEMux
    port map (
            O => \N__33352\,
            I => \N__33338\
        );

    \I__5680\ : Span4Mux_v
    port map (
            O => \N__33349\,
            I => \N__33335\
        );

    \I__5679\ : Span4Mux_v
    port map (
            O => \N__33346\,
            I => \N__33332\
        );

    \I__5678\ : Span4Mux_v
    port map (
            O => \N__33341\,
            I => \N__33329\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__33338\,
            I => \N__33326\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__33335\,
            I => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__5675\ : Odrv4
    port map (
            O => \N__33332\,
            I => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__5674\ : Odrv4
    port map (
            O => \N__33329\,
            I => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__5673\ : Odrv12
    port map (
            O => \N__33326\,
            I => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__5672\ : InMux
    port map (
            O => \N__33317\,
            I => \N__33314\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__33314\,
            I => \phase_controller_inst1.stoper_hc.measured_delay_hc_i_31\
        );

    \I__5670\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33308\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__33308\,
            I => \N__33304\
        );

    \I__5668\ : InMux
    port map (
            O => \N__33307\,
            I => \N__33301\
        );

    \I__5667\ : Span4Mux_h
    port map (
            O => \N__33304\,
            I => \N__33298\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__33301\,
            I => \N__33295\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__33298\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_1
        );

    \I__5664\ : Odrv4
    port map (
            O => \N__33295\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_1
        );

    \I__5663\ : InMux
    port map (
            O => \N__33290\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0\
        );

    \I__5662\ : InMux
    port map (
            O => \N__33287\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1\
        );

    \I__5661\ : InMux
    port map (
            O => \N__33284\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2\
        );

    \I__5660\ : InMux
    port map (
            O => \N__33281\,
            I => \N__33278\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__33278\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_11\
        );

    \I__5658\ : CascadeMux
    port map (
            O => \N__33275\,
            I => \N__33272\
        );

    \I__5657\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33269\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__33269\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_9\
        );

    \I__5655\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33263\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__33263\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_4\
        );

    \I__5653\ : CascadeMux
    port map (
            O => \N__33260\,
            I => \N__33257\
        );

    \I__5652\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33254\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__33254\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_7\
        );

    \I__5650\ : CascadeMux
    port map (
            O => \N__33251\,
            I => \N__33248\
        );

    \I__5649\ : InMux
    port map (
            O => \N__33248\,
            I => \N__33245\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__33245\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_6\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__33242\,
            I => \N__33239\
        );

    \I__5646\ : InMux
    port map (
            O => \N__33239\,
            I => \N__33236\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__33236\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_3\
        );

    \I__5644\ : InMux
    port map (
            O => \N__33233\,
            I => \N__33230\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__33230\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_10\
        );

    \I__5642\ : InMux
    port map (
            O => \N__33227\,
            I => \N__33221\
        );

    \I__5641\ : InMux
    port map (
            O => \N__33226\,
            I => \N__33221\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__33221\,
            I => \N__33218\
        );

    \I__5639\ : Odrv4
    port map (
            O => \N__33218\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_21\
        );

    \I__5638\ : InMux
    port map (
            O => \N__33215\,
            I => \N__33212\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__33212\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_12\
        );

    \I__5636\ : InMux
    port map (
            O => \N__33209\,
            I => \N__33206\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__33206\,
            I => \N__33203\
        );

    \I__5634\ : Span4Mux_v
    port map (
            O => \N__33203\,
            I => \N__33199\
        );

    \I__5633\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33196\
        );

    \I__5632\ : Odrv4
    port map (
            O => \N__33199\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__33196\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__5630\ : InMux
    port map (
            O => \N__33191\,
            I => \bfn_11_23_0_\
        );

    \I__5629\ : InMux
    port map (
            O => \N__33188\,
            I => \N__33185\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__33185\,
            I => \N__33181\
        );

    \I__5627\ : CascadeMux
    port map (
            O => \N__33184\,
            I => \N__33178\
        );

    \I__5626\ : Span4Mux_v
    port map (
            O => \N__33181\,
            I => \N__33175\
        );

    \I__5625\ : InMux
    port map (
            O => \N__33178\,
            I => \N__33172\
        );

    \I__5624\ : Odrv4
    port map (
            O => \N__33175\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__33172\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__5622\ : InMux
    port map (
            O => \N__33167\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__5621\ : InMux
    port map (
            O => \N__33164\,
            I => \N__33161\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__33161\,
            I => \N__33158\
        );

    \I__5619\ : Span4Mux_v
    port map (
            O => \N__33158\,
            I => \N__33154\
        );

    \I__5618\ : InMux
    port map (
            O => \N__33157\,
            I => \N__33151\
        );

    \I__5617\ : Odrv4
    port map (
            O => \N__33154\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__33151\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__5615\ : InMux
    port map (
            O => \N__33146\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__5614\ : InMux
    port map (
            O => \N__33143\,
            I => \N__33140\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__33140\,
            I => \N__33137\
        );

    \I__5612\ : Span4Mux_v
    port map (
            O => \N__33137\,
            I => \N__33134\
        );

    \I__5611\ : Span4Mux_v
    port map (
            O => \N__33134\,
            I => \N__33130\
        );

    \I__5610\ : InMux
    port map (
            O => \N__33133\,
            I => \N__33127\
        );

    \I__5609\ : Odrv4
    port map (
            O => \N__33130\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__33127\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__5607\ : InMux
    port map (
            O => \N__33122\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__5606\ : InMux
    port map (
            O => \N__33119\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__5605\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33113\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__33113\,
            I => \N__33109\
        );

    \I__5603\ : InMux
    port map (
            O => \N__33112\,
            I => \N__33106\
        );

    \I__5602\ : Span4Mux_v
    port map (
            O => \N__33109\,
            I => \N__33103\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__33106\,
            I => \N__33100\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__33103\,
            I => \N__33095\
        );

    \I__5599\ : Span4Mux_v
    port map (
            O => \N__33100\,
            I => \N__33095\
        );

    \I__5598\ : Span4Mux_v
    port map (
            O => \N__33095\,
            I => \N__33092\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__33092\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__5596\ : InMux
    port map (
            O => \N__33089\,
            I => \N__33086\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__33086\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_2\
        );

    \I__5594\ : InMux
    port map (
            O => \N__33083\,
            I => \N__33080\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__33080\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_1\
        );

    \I__5592\ : CascadeMux
    port map (
            O => \N__33077\,
            I => \N__33074\
        );

    \I__5591\ : InMux
    port map (
            O => \N__33074\,
            I => \N__33071\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__33071\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_5\
        );

    \I__5589\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33065\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__33065\,
            I => \N__33062\
        );

    \I__5587\ : Span4Mux_v
    port map (
            O => \N__33062\,
            I => \N__33058\
        );

    \I__5586\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33055\
        );

    \I__5585\ : Odrv4
    port map (
            O => \N__33058\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__33055\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__5583\ : InMux
    port map (
            O => \N__33050\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__5582\ : InMux
    port map (
            O => \N__33047\,
            I => \N__33041\
        );

    \I__5581\ : InMux
    port map (
            O => \N__33046\,
            I => \N__33041\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__33041\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__5579\ : InMux
    port map (
            O => \N__33038\,
            I => \bfn_11_22_0_\
        );

    \I__5578\ : InMux
    port map (
            O => \N__33035\,
            I => \N__33032\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__33032\,
            I => \N__33029\
        );

    \I__5576\ : Span4Mux_h
    port map (
            O => \N__33029\,
            I => \N__33026\
        );

    \I__5575\ : Span4Mux_v
    port map (
            O => \N__33026\,
            I => \N__33022\
        );

    \I__5574\ : InMux
    port map (
            O => \N__33025\,
            I => \N__33019\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__33022\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__33019\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__5571\ : InMux
    port map (
            O => \N__33014\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__5570\ : InMux
    port map (
            O => \N__33011\,
            I => \N__33008\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__33008\,
            I => \N__33005\
        );

    \I__5568\ : Span4Mux_v
    port map (
            O => \N__33005\,
            I => \N__33002\
        );

    \I__5567\ : Span4Mux_v
    port map (
            O => \N__33002\,
            I => \N__32998\
        );

    \I__5566\ : InMux
    port map (
            O => \N__33001\,
            I => \N__32995\
        );

    \I__5565\ : Odrv4
    port map (
            O => \N__32998\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__32995\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__5563\ : InMux
    port map (
            O => \N__32990\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__5562\ : InMux
    port map (
            O => \N__32987\,
            I => \N__32984\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__32984\,
            I => \N__32980\
        );

    \I__5560\ : CascadeMux
    port map (
            O => \N__32983\,
            I => \N__32977\
        );

    \I__5559\ : Span4Mux_v
    port map (
            O => \N__32980\,
            I => \N__32974\
        );

    \I__5558\ : InMux
    port map (
            O => \N__32977\,
            I => \N__32971\
        );

    \I__5557\ : Odrv4
    port map (
            O => \N__32974\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__32971\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__5555\ : InMux
    port map (
            O => \N__32966\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__5554\ : InMux
    port map (
            O => \N__32963\,
            I => \N__32960\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__32960\,
            I => \N__32957\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__32957\,
            I => \N__32954\
        );

    \I__5551\ : Span4Mux_v
    port map (
            O => \N__32954\,
            I => \N__32951\
        );

    \I__5550\ : Span4Mux_v
    port map (
            O => \N__32951\,
            I => \N__32947\
        );

    \I__5549\ : InMux
    port map (
            O => \N__32950\,
            I => \N__32944\
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__32947\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__32944\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__5546\ : InMux
    port map (
            O => \N__32939\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__5545\ : InMux
    port map (
            O => \N__32936\,
            I => \N__32933\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__32933\,
            I => \N__32929\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__32932\,
            I => \N__32926\
        );

    \I__5542\ : Span12Mux_v
    port map (
            O => \N__32929\,
            I => \N__32923\
        );

    \I__5541\ : InMux
    port map (
            O => \N__32926\,
            I => \N__32920\
        );

    \I__5540\ : Odrv12
    port map (
            O => \N__32923\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__32920\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__5538\ : InMux
    port map (
            O => \N__32915\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__5537\ : InMux
    port map (
            O => \N__32912\,
            I => \N__32909\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__32909\,
            I => \N__32906\
        );

    \I__5535\ : Span4Mux_v
    port map (
            O => \N__32906\,
            I => \N__32902\
        );

    \I__5534\ : InMux
    port map (
            O => \N__32905\,
            I => \N__32899\
        );

    \I__5533\ : Odrv4
    port map (
            O => \N__32902\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__32899\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__5531\ : InMux
    port map (
            O => \N__32894\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__5530\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32888\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__32888\,
            I => \N__32885\
        );

    \I__5528\ : Span4Mux_v
    port map (
            O => \N__32885\,
            I => \N__32881\
        );

    \I__5527\ : InMux
    port map (
            O => \N__32884\,
            I => \N__32878\
        );

    \I__5526\ : Odrv4
    port map (
            O => \N__32881\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__32878\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__5524\ : InMux
    port map (
            O => \N__32873\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__5523\ : InMux
    port map (
            O => \N__32870\,
            I => \N__32867\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__32867\,
            I => \N__32864\
        );

    \I__5521\ : Span4Mux_v
    port map (
            O => \N__32864\,
            I => \N__32860\
        );

    \I__5520\ : InMux
    port map (
            O => \N__32863\,
            I => \N__32857\
        );

    \I__5519\ : Odrv4
    port map (
            O => \N__32860\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__32857\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__5517\ : InMux
    port map (
            O => \N__32852\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__5516\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32846\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__32846\,
            I => \N__32843\
        );

    \I__5514\ : Span4Mux_h
    port map (
            O => \N__32843\,
            I => \N__32840\
        );

    \I__5513\ : Span4Mux_v
    port map (
            O => \N__32840\,
            I => \N__32836\
        );

    \I__5512\ : InMux
    port map (
            O => \N__32839\,
            I => \N__32833\
        );

    \I__5511\ : Odrv4
    port map (
            O => \N__32836\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__32833\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__5509\ : InMux
    port map (
            O => \N__32828\,
            I => \bfn_11_21_0_\
        );

    \I__5508\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32822\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__32822\,
            I => \N__32819\
        );

    \I__5506\ : Span4Mux_v
    port map (
            O => \N__32819\,
            I => \N__32815\
        );

    \I__5505\ : InMux
    port map (
            O => \N__32818\,
            I => \N__32812\
        );

    \I__5504\ : Odrv4
    port map (
            O => \N__32815\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__32812\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__5502\ : InMux
    port map (
            O => \N__32807\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__5501\ : InMux
    port map (
            O => \N__32804\,
            I => \N__32801\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__32801\,
            I => \N__32798\
        );

    \I__5499\ : Span4Mux_h
    port map (
            O => \N__32798\,
            I => \N__32795\
        );

    \I__5498\ : Span4Mux_v
    port map (
            O => \N__32795\,
            I => \N__32792\
        );

    \I__5497\ : Span4Mux_v
    port map (
            O => \N__32792\,
            I => \N__32788\
        );

    \I__5496\ : InMux
    port map (
            O => \N__32791\,
            I => \N__32785\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__32788\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__32785\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__5493\ : InMux
    port map (
            O => \N__32780\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__5492\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32774\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__32774\,
            I => \N__32771\
        );

    \I__5490\ : Span4Mux_h
    port map (
            O => \N__32771\,
            I => \N__32768\
        );

    \I__5489\ : Span4Mux_v
    port map (
            O => \N__32768\,
            I => \N__32764\
        );

    \I__5488\ : InMux
    port map (
            O => \N__32767\,
            I => \N__32761\
        );

    \I__5487\ : Odrv4
    port map (
            O => \N__32764\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__32761\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__5485\ : InMux
    port map (
            O => \N__32756\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__5484\ : InMux
    port map (
            O => \N__32753\,
            I => \N__32750\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__32750\,
            I => \N__32747\
        );

    \I__5482\ : Span4Mux_h
    port map (
            O => \N__32747\,
            I => \N__32744\
        );

    \I__5481\ : Span4Mux_v
    port map (
            O => \N__32744\,
            I => \N__32740\
        );

    \I__5480\ : InMux
    port map (
            O => \N__32743\,
            I => \N__32737\
        );

    \I__5479\ : Odrv4
    port map (
            O => \N__32740\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__32737\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__5477\ : InMux
    port map (
            O => \N__32732\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__5476\ : InMux
    port map (
            O => \N__32729\,
            I => \N__32726\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__32726\,
            I => \N__32722\
        );

    \I__5474\ : CascadeMux
    port map (
            O => \N__32725\,
            I => \N__32719\
        );

    \I__5473\ : Span4Mux_v
    port map (
            O => \N__32722\,
            I => \N__32716\
        );

    \I__5472\ : InMux
    port map (
            O => \N__32719\,
            I => \N__32713\
        );

    \I__5471\ : Odrv4
    port map (
            O => \N__32716\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__32713\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__5469\ : InMux
    port map (
            O => \N__32708\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__5468\ : InMux
    port map (
            O => \N__32705\,
            I => \N__32702\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__32702\,
            I => \N__32699\
        );

    \I__5466\ : Span4Mux_v
    port map (
            O => \N__32699\,
            I => \N__32695\
        );

    \I__5465\ : InMux
    port map (
            O => \N__32698\,
            I => \N__32692\
        );

    \I__5464\ : Odrv4
    port map (
            O => \N__32695\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__32692\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__5462\ : InMux
    port map (
            O => \N__32687\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__5461\ : InMux
    port map (
            O => \N__32684\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_29\
        );

    \I__5460\ : InMux
    port map (
            O => \N__32681\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_30\
        );

    \I__5459\ : CEMux
    port map (
            O => \N__32678\,
            I => \N__32672\
        );

    \I__5458\ : CEMux
    port map (
            O => \N__32677\,
            I => \N__32669\
        );

    \I__5457\ : CEMux
    port map (
            O => \N__32676\,
            I => \N__32666\
        );

    \I__5456\ : CEMux
    port map (
            O => \N__32675\,
            I => \N__32663\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__32672\,
            I => \N__32660\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__32669\,
            I => \N__32655\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__32666\,
            I => \N__32655\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__32663\,
            I => \N__32652\
        );

    \I__5451\ : Span4Mux_v
    port map (
            O => \N__32660\,
            I => \N__32647\
        );

    \I__5450\ : Span4Mux_v
    port map (
            O => \N__32655\,
            I => \N__32647\
        );

    \I__5449\ : Span12Mux_h
    port map (
            O => \N__32652\,
            I => \N__32644\
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__32647\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__5447\ : Odrv12
    port map (
            O => \N__32644\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__5446\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32633\
        );

    \I__5445\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32633\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__32633\,
            I => \N__32630\
        );

    \I__5443\ : Span4Mux_h
    port map (
            O => \N__32630\,
            I => \N__32627\
        );

    \I__5442\ : Span4Mux_v
    port map (
            O => \N__32627\,
            I => \N__32624\
        );

    \I__5441\ : Odrv4
    port map (
            O => \N__32624\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__5440\ : CascadeMux
    port map (
            O => \N__32621\,
            I => \N__32618\
        );

    \I__5439\ : InMux
    port map (
            O => \N__32618\,
            I => \N__32614\
        );

    \I__5438\ : InMux
    port map (
            O => \N__32617\,
            I => \N__32611\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__32614\,
            I => \N__32608\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__32611\,
            I => \N__32603\
        );

    \I__5435\ : Span4Mux_h
    port map (
            O => \N__32608\,
            I => \N__32603\
        );

    \I__5434\ : Span4Mux_v
    port map (
            O => \N__32603\,
            I => \N__32600\
        );

    \I__5433\ : Odrv4
    port map (
            O => \N__32600\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__5432\ : InMux
    port map (
            O => \N__32597\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__5431\ : InMux
    port map (
            O => \N__32594\,
            I => \N__32591\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__32591\,
            I => \N__32588\
        );

    \I__5429\ : Span4Mux_v
    port map (
            O => \N__32588\,
            I => \N__32584\
        );

    \I__5428\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32581\
        );

    \I__5427\ : Odrv4
    port map (
            O => \N__32584\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__32581\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__5425\ : InMux
    port map (
            O => \N__32576\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__5424\ : InMux
    port map (
            O => \N__32573\,
            I => \N__32570\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__32570\,
            I => \N__32567\
        );

    \I__5422\ : Span4Mux_v
    port map (
            O => \N__32567\,
            I => \N__32563\
        );

    \I__5421\ : InMux
    port map (
            O => \N__32566\,
            I => \N__32560\
        );

    \I__5420\ : Odrv4
    port map (
            O => \N__32563\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__32560\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__5418\ : InMux
    port map (
            O => \N__32555\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__5417\ : InMux
    port map (
            O => \N__32552\,
            I => \N__32549\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__32549\,
            I => \N__32545\
        );

    \I__5415\ : InMux
    port map (
            O => \N__32548\,
            I => \N__32542\
        );

    \I__5414\ : Span4Mux_h
    port map (
            O => \N__32545\,
            I => \N__32537\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__32542\,
            I => \N__32537\
        );

    \I__5412\ : Span4Mux_v
    port map (
            O => \N__32537\,
            I => \N__32534\
        );

    \I__5411\ : Odrv4
    port map (
            O => \N__32534\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__5410\ : InMux
    port map (
            O => \N__32531\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__32528\,
            I => \N__32524\
        );

    \I__5408\ : InMux
    port map (
            O => \N__32527\,
            I => \N__32519\
        );

    \I__5407\ : InMux
    port map (
            O => \N__32524\,
            I => \N__32519\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__32519\,
            I => \N__32516\
        );

    \I__5405\ : Span12Mux_v
    port map (
            O => \N__32516\,
            I => \N__32513\
        );

    \I__5404\ : Odrv12
    port map (
            O => \N__32513\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__5403\ : InMux
    port map (
            O => \N__32510\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__5402\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32504\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__32504\,
            I => \N__32500\
        );

    \I__5400\ : CascadeMux
    port map (
            O => \N__32503\,
            I => \N__32497\
        );

    \I__5399\ : Span4Mux_v
    port map (
            O => \N__32500\,
            I => \N__32494\
        );

    \I__5398\ : InMux
    port map (
            O => \N__32497\,
            I => \N__32491\
        );

    \I__5397\ : Odrv4
    port map (
            O => \N__32494\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__32491\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__5395\ : InMux
    port map (
            O => \N__32486\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__5394\ : CascadeMux
    port map (
            O => \N__32483\,
            I => \N__32479\
        );

    \I__5393\ : CascadeMux
    port map (
            O => \N__32482\,
            I => \N__32476\
        );

    \I__5392\ : InMux
    port map (
            O => \N__32479\,
            I => \N__32471\
        );

    \I__5391\ : InMux
    port map (
            O => \N__32476\,
            I => \N__32471\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__32471\,
            I => \N__32467\
        );

    \I__5389\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32464\
        );

    \I__5388\ : Span12Mux_s11_v
    port map (
            O => \N__32467\,
            I => \N__32461\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__32464\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_22\
        );

    \I__5386\ : Odrv12
    port map (
            O => \N__32461\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_22\
        );

    \I__5385\ : InMux
    port map (
            O => \N__32456\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_21\
        );

    \I__5384\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32447\
        );

    \I__5383\ : InMux
    port map (
            O => \N__32452\,
            I => \N__32447\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__32447\,
            I => \N__32443\
        );

    \I__5381\ : InMux
    port map (
            O => \N__32446\,
            I => \N__32440\
        );

    \I__5380\ : Span12Mux_v
    port map (
            O => \N__32443\,
            I => \N__32437\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__32440\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_23\
        );

    \I__5378\ : Odrv12
    port map (
            O => \N__32437\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_23\
        );

    \I__5377\ : InMux
    port map (
            O => \N__32432\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_22\
        );

    \I__5376\ : CascadeMux
    port map (
            O => \N__32429\,
            I => \N__32425\
        );

    \I__5375\ : CascadeMux
    port map (
            O => \N__32428\,
            I => \N__32422\
        );

    \I__5374\ : InMux
    port map (
            O => \N__32425\,
            I => \N__32417\
        );

    \I__5373\ : InMux
    port map (
            O => \N__32422\,
            I => \N__32417\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__32417\,
            I => \N__32413\
        );

    \I__5371\ : InMux
    port map (
            O => \N__32416\,
            I => \N__32410\
        );

    \I__5370\ : Span12Mux_v
    port map (
            O => \N__32413\,
            I => \N__32407\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__32410\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_24\
        );

    \I__5368\ : Odrv12
    port map (
            O => \N__32407\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_24\
        );

    \I__5367\ : InMux
    port map (
            O => \N__32402\,
            I => \bfn_11_19_0_\
        );

    \I__5366\ : InMux
    port map (
            O => \N__32399\,
            I => \N__32393\
        );

    \I__5365\ : InMux
    port map (
            O => \N__32398\,
            I => \N__32393\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__32393\,
            I => \N__32389\
        );

    \I__5363\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32386\
        );

    \I__5362\ : Span12Mux_v
    port map (
            O => \N__32389\,
            I => \N__32383\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__32386\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_25\
        );

    \I__5360\ : Odrv12
    port map (
            O => \N__32383\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_25\
        );

    \I__5359\ : InMux
    port map (
            O => \N__32378\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_24\
        );

    \I__5358\ : CascadeMux
    port map (
            O => \N__32375\,
            I => \N__32371\
        );

    \I__5357\ : CascadeMux
    port map (
            O => \N__32374\,
            I => \N__32368\
        );

    \I__5356\ : InMux
    port map (
            O => \N__32371\,
            I => \N__32362\
        );

    \I__5355\ : InMux
    port map (
            O => \N__32368\,
            I => \N__32362\
        );

    \I__5354\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32359\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__32362\,
            I => \N__32356\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__32359\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_26\
        );

    \I__5351\ : Odrv12
    port map (
            O => \N__32356\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_26\
        );

    \I__5350\ : InMux
    port map (
            O => \N__32351\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_25\
        );

    \I__5349\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32341\
        );

    \I__5348\ : InMux
    port map (
            O => \N__32347\,
            I => \N__32341\
        );

    \I__5347\ : InMux
    port map (
            O => \N__32346\,
            I => \N__32338\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__32341\,
            I => \N__32335\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__32338\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_27\
        );

    \I__5344\ : Odrv12
    port map (
            O => \N__32335\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_27\
        );

    \I__5343\ : InMux
    port map (
            O => \N__32330\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_26\
        );

    \I__5342\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32321\
        );

    \I__5341\ : InMux
    port map (
            O => \N__32326\,
            I => \N__32321\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__32321\,
            I => \N__32317\
        );

    \I__5339\ : InMux
    port map (
            O => \N__32320\,
            I => \N__32314\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__32317\,
            I => \N__32311\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__32314\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_28\
        );

    \I__5336\ : Odrv4
    port map (
            O => \N__32311\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_28\
        );

    \I__5335\ : InMux
    port map (
            O => \N__32306\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_27\
        );

    \I__5334\ : InMux
    port map (
            O => \N__32303\,
            I => \N__32297\
        );

    \I__5333\ : InMux
    port map (
            O => \N__32302\,
            I => \N__32297\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__32297\,
            I => \N__32293\
        );

    \I__5331\ : InMux
    port map (
            O => \N__32296\,
            I => \N__32290\
        );

    \I__5330\ : Span4Mux_v
    port map (
            O => \N__32293\,
            I => \N__32287\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__32290\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_29\
        );

    \I__5328\ : Odrv4
    port map (
            O => \N__32287\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_29\
        );

    \I__5327\ : InMux
    port map (
            O => \N__32282\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_28\
        );

    \I__5326\ : InMux
    port map (
            O => \N__32279\,
            I => \N__32276\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__32276\,
            I => \N__32272\
        );

    \I__5324\ : InMux
    port map (
            O => \N__32275\,
            I => \N__32269\
        );

    \I__5323\ : Span4Mux_v
    port map (
            O => \N__32272\,
            I => \N__32266\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__32269\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_13\
        );

    \I__5321\ : Odrv4
    port map (
            O => \N__32266\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_13\
        );

    \I__5320\ : InMux
    port map (
            O => \N__32261\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_12\
        );

    \I__5319\ : InMux
    port map (
            O => \N__32258\,
            I => \N__32254\
        );

    \I__5318\ : InMux
    port map (
            O => \N__32257\,
            I => \N__32251\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__32254\,
            I => \N__32248\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__32251\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_14\
        );

    \I__5315\ : Odrv12
    port map (
            O => \N__32248\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_14\
        );

    \I__5314\ : InMux
    port map (
            O => \N__32243\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_13\
        );

    \I__5313\ : InMux
    port map (
            O => \N__32240\,
            I => \N__32236\
        );

    \I__5312\ : InMux
    port map (
            O => \N__32239\,
            I => \N__32233\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__32236\,
            I => \N__32230\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__32233\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_15\
        );

    \I__5309\ : Odrv12
    port map (
            O => \N__32230\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_15\
        );

    \I__5308\ : InMux
    port map (
            O => \N__32225\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_14\
        );

    \I__5307\ : InMux
    port map (
            O => \N__32222\,
            I => \bfn_11_18_0_\
        );

    \I__5306\ : InMux
    port map (
            O => \N__32219\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_16\
        );

    \I__5305\ : InMux
    port map (
            O => \N__32216\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_17\
        );

    \I__5304\ : InMux
    port map (
            O => \N__32213\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_18\
        );

    \I__5303\ : CascadeMux
    port map (
            O => \N__32210\,
            I => \N__32206\
        );

    \I__5302\ : CascadeMux
    port map (
            O => \N__32209\,
            I => \N__32203\
        );

    \I__5301\ : InMux
    port map (
            O => \N__32206\,
            I => \N__32198\
        );

    \I__5300\ : InMux
    port map (
            O => \N__32203\,
            I => \N__32198\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__32198\,
            I => \N__32194\
        );

    \I__5298\ : InMux
    port map (
            O => \N__32197\,
            I => \N__32191\
        );

    \I__5297\ : Sp12to4
    port map (
            O => \N__32194\,
            I => \N__32188\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__32191\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_20\
        );

    \I__5295\ : Odrv12
    port map (
            O => \N__32188\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_20\
        );

    \I__5294\ : InMux
    port map (
            O => \N__32183\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_19\
        );

    \I__5293\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32174\
        );

    \I__5292\ : InMux
    port map (
            O => \N__32179\,
            I => \N__32174\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__32174\,
            I => \N__32171\
        );

    \I__5290\ : Span4Mux_h
    port map (
            O => \N__32171\,
            I => \N__32167\
        );

    \I__5289\ : InMux
    port map (
            O => \N__32170\,
            I => \N__32164\
        );

    \I__5288\ : Span4Mux_v
    port map (
            O => \N__32167\,
            I => \N__32161\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__32164\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_21\
        );

    \I__5286\ : Odrv4
    port map (
            O => \N__32161\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_21\
        );

    \I__5285\ : InMux
    port map (
            O => \N__32156\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_20\
        );

    \I__5284\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32149\
        );

    \I__5283\ : InMux
    port map (
            O => \N__32152\,
            I => \N__32146\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__32149\,
            I => \N__32143\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__32146\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_5\
        );

    \I__5280\ : Odrv12
    port map (
            O => \N__32143\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_5\
        );

    \I__5279\ : InMux
    port map (
            O => \N__32138\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_4\
        );

    \I__5278\ : InMux
    port map (
            O => \N__32135\,
            I => \N__32132\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__32132\,
            I => \N__32128\
        );

    \I__5276\ : InMux
    port map (
            O => \N__32131\,
            I => \N__32125\
        );

    \I__5275\ : Span4Mux_v
    port map (
            O => \N__32128\,
            I => \N__32122\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__32125\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_6\
        );

    \I__5273\ : Odrv4
    port map (
            O => \N__32122\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_6\
        );

    \I__5272\ : InMux
    port map (
            O => \N__32117\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_5\
        );

    \I__5271\ : InMux
    port map (
            O => \N__32114\,
            I => \N__32110\
        );

    \I__5270\ : InMux
    port map (
            O => \N__32113\,
            I => \N__32107\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__32110\,
            I => \N__32104\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__32107\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_7\
        );

    \I__5267\ : Odrv12
    port map (
            O => \N__32104\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_7\
        );

    \I__5266\ : InMux
    port map (
            O => \N__32099\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_6\
        );

    \I__5265\ : InMux
    port map (
            O => \N__32096\,
            I => \N__32092\
        );

    \I__5264\ : InMux
    port map (
            O => \N__32095\,
            I => \N__32089\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__32092\,
            I => \N__32086\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__32089\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_8\
        );

    \I__5261\ : Odrv12
    port map (
            O => \N__32086\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_8\
        );

    \I__5260\ : InMux
    port map (
            O => \N__32081\,
            I => \bfn_11_17_0_\
        );

    \I__5259\ : InMux
    port map (
            O => \N__32078\,
            I => \N__32074\
        );

    \I__5258\ : InMux
    port map (
            O => \N__32077\,
            I => \N__32071\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__32074\,
            I => \N__32068\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__32071\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_9\
        );

    \I__5255\ : Odrv12
    port map (
            O => \N__32068\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_9\
        );

    \I__5254\ : InMux
    port map (
            O => \N__32063\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_8\
        );

    \I__5253\ : InMux
    port map (
            O => \N__32060\,
            I => \N__32057\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__32057\,
            I => \N__32053\
        );

    \I__5251\ : InMux
    port map (
            O => \N__32056\,
            I => \N__32050\
        );

    \I__5250\ : Span4Mux_h
    port map (
            O => \N__32053\,
            I => \N__32047\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__32050\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_10\
        );

    \I__5248\ : Odrv4
    port map (
            O => \N__32047\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_10\
        );

    \I__5247\ : InMux
    port map (
            O => \N__32042\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_9\
        );

    \I__5246\ : InMux
    port map (
            O => \N__32039\,
            I => \N__32035\
        );

    \I__5245\ : InMux
    port map (
            O => \N__32038\,
            I => \N__32032\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__32035\,
            I => \N__32029\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__32032\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_11\
        );

    \I__5242\ : Odrv12
    port map (
            O => \N__32029\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_11\
        );

    \I__5241\ : InMux
    port map (
            O => \N__32024\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_10\
        );

    \I__5240\ : InMux
    port map (
            O => \N__32021\,
            I => \N__32018\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__32018\,
            I => \N__32014\
        );

    \I__5238\ : InMux
    port map (
            O => \N__32017\,
            I => \N__32011\
        );

    \I__5237\ : Span4Mux_h
    port map (
            O => \N__32014\,
            I => \N__32008\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__32011\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_12\
        );

    \I__5235\ : Odrv4
    port map (
            O => \N__32008\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_12\
        );

    \I__5234\ : InMux
    port map (
            O => \N__32003\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_11\
        );

    \I__5233\ : CascadeMux
    port map (
            O => \N__32000\,
            I => \N__31997\
        );

    \I__5232\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31994\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__31994\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28\
        );

    \I__5230\ : InMux
    port map (
            O => \N__31991\,
            I => \N__31988\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__31988\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30\
        );

    \I__5228\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31982\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__31982\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt28\
        );

    \I__5226\ : CascadeMux
    port map (
            O => \N__31979\,
            I => \N__31975\
        );

    \I__5225\ : InMux
    port map (
            O => \N__31978\,
            I => \N__31972\
        );

    \I__5224\ : InMux
    port map (
            O => \N__31975\,
            I => \N__31969\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__31972\,
            I => \phase_controller_inst1.stoper_hc.counter\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__31969\,
            I => \phase_controller_inst1.stoper_hc.counter\
        );

    \I__5221\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31961\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__31961\,
            I => \N__31957\
        );

    \I__5219\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31954\
        );

    \I__5218\ : Span4Mux_v
    port map (
            O => \N__31957\,
            I => \N__31951\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__31954\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_0\
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__31951\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_0\
        );

    \I__5215\ : InMux
    port map (
            O => \N__31946\,
            I => \N__31943\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__31943\,
            I => \N__31939\
        );

    \I__5213\ : InMux
    port map (
            O => \N__31942\,
            I => \N__31936\
        );

    \I__5212\ : Span4Mux_v
    port map (
            O => \N__31939\,
            I => \N__31933\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__31936\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_1\
        );

    \I__5210\ : Odrv4
    port map (
            O => \N__31933\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_1\
        );

    \I__5209\ : InMux
    port map (
            O => \N__31928\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_0\
        );

    \I__5208\ : InMux
    port map (
            O => \N__31925\,
            I => \N__31922\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__31922\,
            I => \N__31918\
        );

    \I__5206\ : InMux
    port map (
            O => \N__31921\,
            I => \N__31915\
        );

    \I__5205\ : Span4Mux_v
    port map (
            O => \N__31918\,
            I => \N__31912\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__31915\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_2\
        );

    \I__5203\ : Odrv4
    port map (
            O => \N__31912\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_2\
        );

    \I__5202\ : InMux
    port map (
            O => \N__31907\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_1\
        );

    \I__5201\ : InMux
    port map (
            O => \N__31904\,
            I => \N__31900\
        );

    \I__5200\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31897\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__31900\,
            I => \N__31894\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__31897\,
            I => \N__31889\
        );

    \I__5197\ : Span4Mux_v
    port map (
            O => \N__31894\,
            I => \N__31889\
        );

    \I__5196\ : Odrv4
    port map (
            O => \N__31889\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_3\
        );

    \I__5195\ : InMux
    port map (
            O => \N__31886\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_2\
        );

    \I__5194\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31880\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__31880\,
            I => \N__31876\
        );

    \I__5192\ : InMux
    port map (
            O => \N__31879\,
            I => \N__31873\
        );

    \I__5191\ : Span4Mux_v
    port map (
            O => \N__31876\,
            I => \N__31870\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__31873\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_4\
        );

    \I__5189\ : Odrv4
    port map (
            O => \N__31870\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_4\
        );

    \I__5188\ : InMux
    port map (
            O => \N__31865\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_3\
        );

    \I__5187\ : InMux
    port map (
            O => \N__31862\,
            I => \N__31859\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__31859\,
            I => \N__31856\
        );

    \I__5185\ : Span4Mux_v
    port map (
            O => \N__31856\,
            I => \N__31853\
        );

    \I__5184\ : Odrv4
    port map (
            O => \N__31853\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt22\
        );

    \I__5183\ : CascadeMux
    port map (
            O => \N__31850\,
            I => \N__31847\
        );

    \I__5182\ : InMux
    port map (
            O => \N__31847\,
            I => \N__31844\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__31844\,
            I => \N__31841\
        );

    \I__5180\ : Span4Mux_v
    port map (
            O => \N__31841\,
            I => \N__31838\
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__31838\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22\
        );

    \I__5178\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31832\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__31832\,
            I => \N__31829\
        );

    \I__5176\ : Odrv4
    port map (
            O => \N__31829\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24\
        );

    \I__5175\ : CascadeMux
    port map (
            O => \N__31826\,
            I => \N__31823\
        );

    \I__5174\ : InMux
    port map (
            O => \N__31823\,
            I => \N__31820\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__31820\,
            I => \N__31817\
        );

    \I__5172\ : Odrv12
    port map (
            O => \N__31817\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt24\
        );

    \I__5171\ : InMux
    port map (
            O => \N__31814\,
            I => \N__31811\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__31811\,
            I => \N__31808\
        );

    \I__5169\ : Span4Mux_h
    port map (
            O => \N__31808\,
            I => \N__31805\
        );

    \I__5168\ : Odrv4
    port map (
            O => \N__31805\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt26\
        );

    \I__5167\ : CascadeMux
    port map (
            O => \N__31802\,
            I => \N__31799\
        );

    \I__5166\ : InMux
    port map (
            O => \N__31799\,
            I => \N__31796\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__31796\,
            I => \N__31793\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__31793\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26\
        );

    \I__5163\ : InMux
    port map (
            O => \N__31790\,
            I => \bfn_11_15_0_\
        );

    \I__5162\ : InMux
    port map (
            O => \N__31787\,
            I => \N__31782\
        );

    \I__5161\ : InMux
    port map (
            O => \N__31786\,
            I => \N__31775\
        );

    \I__5160\ : InMux
    port map (
            O => \N__31785\,
            I => \N__31763\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__31782\,
            I => \N__31760\
        );

    \I__5158\ : InMux
    port map (
            O => \N__31781\,
            I => \N__31747\
        );

    \I__5157\ : InMux
    port map (
            O => \N__31780\,
            I => \N__31747\
        );

    \I__5156\ : InMux
    port map (
            O => \N__31779\,
            I => \N__31747\
        );

    \I__5155\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31747\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__31775\,
            I => \N__31744\
        );

    \I__5153\ : InMux
    port map (
            O => \N__31774\,
            I => \N__31737\
        );

    \I__5152\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31737\
        );

    \I__5151\ : InMux
    port map (
            O => \N__31772\,
            I => \N__31737\
        );

    \I__5150\ : InMux
    port map (
            O => \N__31771\,
            I => \N__31720\
        );

    \I__5149\ : InMux
    port map (
            O => \N__31770\,
            I => \N__31720\
        );

    \I__5148\ : InMux
    port map (
            O => \N__31769\,
            I => \N__31720\
        );

    \I__5147\ : InMux
    port map (
            O => \N__31768\,
            I => \N__31713\
        );

    \I__5146\ : InMux
    port map (
            O => \N__31767\,
            I => \N__31713\
        );

    \I__5145\ : InMux
    port map (
            O => \N__31766\,
            I => \N__31713\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__31763\,
            I => \N__31710\
        );

    \I__5143\ : Span4Mux_h
    port map (
            O => \N__31760\,
            I => \N__31707\
        );

    \I__5142\ : InMux
    port map (
            O => \N__31759\,
            I => \N__31698\
        );

    \I__5141\ : InMux
    port map (
            O => \N__31758\,
            I => \N__31698\
        );

    \I__5140\ : InMux
    port map (
            O => \N__31757\,
            I => \N__31698\
        );

    \I__5139\ : InMux
    port map (
            O => \N__31756\,
            I => \N__31698\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__31747\,
            I => \N__31693\
        );

    \I__5137\ : Span12Mux_v
    port map (
            O => \N__31744\,
            I => \N__31693\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__31737\,
            I => \N__31690\
        );

    \I__5135\ : InMux
    port map (
            O => \N__31736\,
            I => \N__31685\
        );

    \I__5134\ : InMux
    port map (
            O => \N__31735\,
            I => \N__31685\
        );

    \I__5133\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31682\
        );

    \I__5132\ : InMux
    port map (
            O => \N__31733\,
            I => \N__31677\
        );

    \I__5131\ : InMux
    port map (
            O => \N__31732\,
            I => \N__31677\
        );

    \I__5130\ : InMux
    port map (
            O => \N__31731\,
            I => \N__31668\
        );

    \I__5129\ : InMux
    port map (
            O => \N__31730\,
            I => \N__31668\
        );

    \I__5128\ : InMux
    port map (
            O => \N__31729\,
            I => \N__31668\
        );

    \I__5127\ : InMux
    port map (
            O => \N__31728\,
            I => \N__31668\
        );

    \I__5126\ : InMux
    port map (
            O => \N__31727\,
            I => \N__31665\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__31720\,
            I => \N__31660\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__31713\,
            I => \N__31660\
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__31710\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__31707\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__31698\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5120\ : Odrv12
    port map (
            O => \N__31693\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5119\ : Odrv4
    port map (
            O => \N__31690\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__31685\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__31682\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__31677\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__31668\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__31665\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5113\ : Odrv4
    port map (
            O => \N__31660\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5112\ : InMux
    port map (
            O => \N__31637\,
            I => \N__31634\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__31634\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__5110\ : CascadeMux
    port map (
            O => \N__31631\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\
        );

    \I__5109\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31625\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__31625\,
            I => \N__31622\
        );

    \I__5107\ : Span4Mux_h
    port map (
            O => \N__31622\,
            I => \N__31619\
        );

    \I__5106\ : Odrv4
    port map (
            O => \N__31619\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22\
        );

    \I__5105\ : CascadeMux
    port map (
            O => \N__31616\,
            I => \N__31613\
        );

    \I__5104\ : InMux
    port map (
            O => \N__31613\,
            I => \N__31610\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__31610\,
            I => \N__31607\
        );

    \I__5102\ : Span4Mux_v
    port map (
            O => \N__31607\,
            I => \N__31604\
        );

    \I__5101\ : Span4Mux_v
    port map (
            O => \N__31604\,
            I => \N__31601\
        );

    \I__5100\ : Odrv4
    port map (
            O => \N__31601\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_11\
        );

    \I__5099\ : InMux
    port map (
            O => \N__31598\,
            I => \N__31595\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__31595\,
            I => \phase_controller_inst1.stoper_hc.counter_i_11\
        );

    \I__5097\ : InMux
    port map (
            O => \N__31592\,
            I => \N__31589\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__31589\,
            I => \N__31586\
        );

    \I__5095\ : Span4Mux_v
    port map (
            O => \N__31586\,
            I => \N__31583\
        );

    \I__5094\ : Odrv4
    port map (
            O => \N__31583\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_12\
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__31580\,
            I => \N__31577\
        );

    \I__5092\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31574\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__31574\,
            I => \phase_controller_inst1.stoper_hc.counter_i_12\
        );

    \I__5090\ : InMux
    port map (
            O => \N__31571\,
            I => \N__31568\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__31568\,
            I => \N__31565\
        );

    \I__5088\ : Odrv12
    port map (
            O => \N__31565\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_13\
        );

    \I__5087\ : CascadeMux
    port map (
            O => \N__31562\,
            I => \N__31559\
        );

    \I__5086\ : InMux
    port map (
            O => \N__31559\,
            I => \N__31556\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__31556\,
            I => \N__31553\
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__31553\,
            I => \phase_controller_inst1.stoper_hc.counter_i_13\
        );

    \I__5083\ : InMux
    port map (
            O => \N__31550\,
            I => \N__31547\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__31547\,
            I => \N__31544\
        );

    \I__5081\ : Span4Mux_v
    port map (
            O => \N__31544\,
            I => \N__31541\
        );

    \I__5080\ : Odrv4
    port map (
            O => \N__31541\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_14\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__31538\,
            I => \N__31535\
        );

    \I__5078\ : InMux
    port map (
            O => \N__31535\,
            I => \N__31532\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__31532\,
            I => \N__31529\
        );

    \I__5076\ : Odrv4
    port map (
            O => \N__31529\,
            I => \phase_controller_inst1.stoper_hc.counter_i_14\
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__31526\,
            I => \N__31523\
        );

    \I__5074\ : InMux
    port map (
            O => \N__31523\,
            I => \N__31520\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__31520\,
            I => \N__31517\
        );

    \I__5072\ : Odrv12
    port map (
            O => \N__31517\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_15\
        );

    \I__5071\ : InMux
    port map (
            O => \N__31514\,
            I => \N__31511\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__31511\,
            I => \phase_controller_inst1.stoper_hc.counter_i_15\
        );

    \I__5069\ : InMux
    port map (
            O => \N__31508\,
            I => \N__31505\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__31505\,
            I => \N__31502\
        );

    \I__5067\ : Odrv12
    port map (
            O => \N__31502\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20\
        );

    \I__5066\ : CascadeMux
    port map (
            O => \N__31499\,
            I => \N__31496\
        );

    \I__5065\ : InMux
    port map (
            O => \N__31496\,
            I => \N__31493\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__31493\,
            I => \N__31490\
        );

    \I__5063\ : Odrv12
    port map (
            O => \N__31490\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt20\
        );

    \I__5062\ : CascadeMux
    port map (
            O => \N__31487\,
            I => \N__31484\
        );

    \I__5061\ : InMux
    port map (
            O => \N__31484\,
            I => \N__31481\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__31481\,
            I => \N__31478\
        );

    \I__5059\ : Odrv4
    port map (
            O => \N__31478\,
            I => \phase_controller_inst1.stoper_hc.counter_i_3\
        );

    \I__5058\ : CascadeMux
    port map (
            O => \N__31475\,
            I => \N__31472\
        );

    \I__5057\ : InMux
    port map (
            O => \N__31472\,
            I => \N__31469\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__31469\,
            I => \N__31466\
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__31466\,
            I => \phase_controller_inst1.stoper_hc.counter_i_4\
        );

    \I__5054\ : InMux
    port map (
            O => \N__31463\,
            I => \N__31460\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__31460\,
            I => \N__31457\
        );

    \I__5052\ : Span4Mux_v
    port map (
            O => \N__31457\,
            I => \N__31454\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__31454\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_5\
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__31451\,
            I => \N__31448\
        );

    \I__5049\ : InMux
    port map (
            O => \N__31448\,
            I => \N__31445\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__31445\,
            I => \N__31442\
        );

    \I__5047\ : Odrv12
    port map (
            O => \N__31442\,
            I => \phase_controller_inst1.stoper_hc.counter_i_5\
        );

    \I__5046\ : InMux
    port map (
            O => \N__31439\,
            I => \N__31436\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__31436\,
            I => \phase_controller_inst1.stoper_hc.counter_i_6\
        );

    \I__5044\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31430\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__31430\,
            I => \phase_controller_inst1.stoper_hc.counter_i_7\
        );

    \I__5042\ : InMux
    port map (
            O => \N__31427\,
            I => \N__31424\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__31424\,
            I => \N__31421\
        );

    \I__5040\ : Odrv12
    port map (
            O => \N__31421\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_8\
        );

    \I__5039\ : CascadeMux
    port map (
            O => \N__31418\,
            I => \N__31415\
        );

    \I__5038\ : InMux
    port map (
            O => \N__31415\,
            I => \N__31412\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__31412\,
            I => \phase_controller_inst1.stoper_hc.counter_i_8\
        );

    \I__5036\ : InMux
    port map (
            O => \N__31409\,
            I => \N__31406\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__31406\,
            I => \N__31403\
        );

    \I__5034\ : Odrv12
    port map (
            O => \N__31403\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_9\
        );

    \I__5033\ : CascadeMux
    port map (
            O => \N__31400\,
            I => \N__31397\
        );

    \I__5032\ : InMux
    port map (
            O => \N__31397\,
            I => \N__31394\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__31394\,
            I => \phase_controller_inst1.stoper_hc.counter_i_9\
        );

    \I__5030\ : CascadeMux
    port map (
            O => \N__31391\,
            I => \N__31388\
        );

    \I__5029\ : InMux
    port map (
            O => \N__31388\,
            I => \N__31385\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__31385\,
            I => \phase_controller_inst1.stoper_hc.counter_i_10\
        );

    \I__5027\ : InMux
    port map (
            O => \N__31382\,
            I => \N__31376\
        );

    \I__5026\ : InMux
    port map (
            O => \N__31381\,
            I => \N__31376\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__31376\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24\
        );

    \I__5024\ : InMux
    port map (
            O => \N__31373\,
            I => \N__31367\
        );

    \I__5023\ : InMux
    port map (
            O => \N__31372\,
            I => \N__31367\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__31367\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_26\
        );

    \I__5021\ : InMux
    port map (
            O => \N__31364\,
            I => \N__31358\
        );

    \I__5020\ : InMux
    port map (
            O => \N__31363\,
            I => \N__31358\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__31358\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_27\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__31355\,
            I => \N__31352\
        );

    \I__5017\ : InMux
    port map (
            O => \N__31352\,
            I => \N__31349\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__31349\,
            I => \phase_controller_inst1.stoper_hc.counter_i_0\
        );

    \I__5015\ : CascadeMux
    port map (
            O => \N__31346\,
            I => \N__31343\
        );

    \I__5014\ : InMux
    port map (
            O => \N__31343\,
            I => \N__31340\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__31340\,
            I => \N__31337\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__31337\,
            I => \N__31334\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__31334\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ1Z_1\
        );

    \I__5010\ : InMux
    port map (
            O => \N__31331\,
            I => \N__31328\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__31328\,
            I => \phase_controller_inst1.stoper_hc.counter_i_1\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__31325\,
            I => \N__31322\
        );

    \I__5007\ : InMux
    port map (
            O => \N__31322\,
            I => \N__31319\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__31319\,
            I => \phase_controller_inst1.stoper_hc.counter_i_2\
        );

    \I__5005\ : InMux
    port map (
            O => \N__31316\,
            I => \N__31310\
        );

    \I__5004\ : InMux
    port map (
            O => \N__31315\,
            I => \N__31310\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__31310\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_17\
        );

    \I__5002\ : InMux
    port map (
            O => \N__31307\,
            I => \N__31301\
        );

    \I__5001\ : InMux
    port map (
            O => \N__31306\,
            I => \N__31301\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__31301\,
            I => \N__31298\
        );

    \I__4999\ : Odrv4
    port map (
            O => \N__31298\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_24\
        );

    \I__4998\ : InMux
    port map (
            O => \N__31295\,
            I => \N__31289\
        );

    \I__4997\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31289\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__31289\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_20\
        );

    \I__4995\ : InMux
    port map (
            O => \N__31286\,
            I => \N__31280\
        );

    \I__4994\ : InMux
    port map (
            O => \N__31285\,
            I => \N__31280\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__31280\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_21\
        );

    \I__4992\ : InMux
    port map (
            O => \N__31277\,
            I => \N__31271\
        );

    \I__4991\ : InMux
    port map (
            O => \N__31276\,
            I => \N__31271\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__31271\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_22\
        );

    \I__4989\ : InMux
    port map (
            O => \N__31268\,
            I => \N__31262\
        );

    \I__4988\ : InMux
    port map (
            O => \N__31267\,
            I => \N__31262\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__31262\,
            I => \N__31259\
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__31259\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_23\
        );

    \I__4985\ : InMux
    port map (
            O => \N__31256\,
            I => \N__31250\
        );

    \I__4984\ : InMux
    port map (
            O => \N__31255\,
            I => \N__31250\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__31250\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_23\
        );

    \I__4982\ : InMux
    port map (
            O => \N__31247\,
            I => \N__31241\
        );

    \I__4981\ : InMux
    port map (
            O => \N__31246\,
            I => \N__31241\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__31241\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_22\
        );

    \I__4979\ : InMux
    port map (
            O => \N__31238\,
            I => \N__31235\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__31235\,
            I => \N__31231\
        );

    \I__4977\ : InMux
    port map (
            O => \N__31234\,
            I => \N__31228\
        );

    \I__4976\ : Span4Mux_h
    port map (
            O => \N__31231\,
            I => \N__31225\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__31228\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19\
        );

    \I__4974\ : Odrv4
    port map (
            O => \N__31225\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19\
        );

    \I__4973\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31214\
        );

    \I__4972\ : InMux
    port map (
            O => \N__31219\,
            I => \N__31214\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__31214\,
            I => \N__31211\
        );

    \I__4970\ : Odrv4
    port map (
            O => \N__31211\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_20\
        );

    \I__4969\ : CascadeMux
    port map (
            O => \N__31208\,
            I => \N__31204\
        );

    \I__4968\ : CascadeMux
    port map (
            O => \N__31207\,
            I => \N__31201\
        );

    \I__4967\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31196\
        );

    \I__4966\ : InMux
    port map (
            O => \N__31201\,
            I => \N__31196\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__31196\,
            I => \N__31193\
        );

    \I__4964\ : Odrv4
    port map (
            O => \N__31193\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_25\
        );

    \I__4963\ : CascadeMux
    port map (
            O => \N__31190\,
            I => \N__31186\
        );

    \I__4962\ : CascadeMux
    port map (
            O => \N__31189\,
            I => \N__31183\
        );

    \I__4961\ : InMux
    port map (
            O => \N__31186\,
            I => \N__31178\
        );

    \I__4960\ : InMux
    port map (
            O => \N__31183\,
            I => \N__31178\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__31178\,
            I => \N__31175\
        );

    \I__4958\ : Odrv4
    port map (
            O => \N__31175\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_27\
        );

    \I__4957\ : InMux
    port map (
            O => \N__31172\,
            I => \N__31169\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__31169\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__31166\,
            I => \N__31163\
        );

    \I__4954\ : InMux
    port map (
            O => \N__31163\,
            I => \N__31160\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__31160\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt26\
        );

    \I__4952\ : InMux
    port map (
            O => \N__31157\,
            I => \N__31154\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__31154\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt28\
        );

    \I__4950\ : CascadeMux
    port map (
            O => \N__31151\,
            I => \N__31148\
        );

    \I__4949\ : InMux
    port map (
            O => \N__31148\,
            I => \N__31145\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__31145\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28\
        );

    \I__4947\ : InMux
    port map (
            O => \N__31142\,
            I => \N__31139\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__31139\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt30\
        );

    \I__4945\ : CascadeMux
    port map (
            O => \N__31136\,
            I => \N__31133\
        );

    \I__4944\ : InMux
    port map (
            O => \N__31133\,
            I => \N__31130\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__31130\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30\
        );

    \I__4942\ : InMux
    port map (
            O => \N__31127\,
            I => \bfn_11_7_0_\
        );

    \I__4941\ : CascadeMux
    port map (
            O => \N__31124\,
            I => \N__31119\
        );

    \I__4940\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31116\
        );

    \I__4939\ : InMux
    port map (
            O => \N__31122\,
            I => \N__31111\
        );

    \I__4938\ : InMux
    port map (
            O => \N__31119\,
            I => \N__31111\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__31116\,
            I => \N__31108\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__31111\,
            I => \N__31105\
        );

    \I__4935\ : Span4Mux_s2_v
    port map (
            O => \N__31108\,
            I => \N__31102\
        );

    \I__4934\ : Odrv4
    port map (
            O => \N__31105\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\
        );

    \I__4933\ : Odrv4
    port map (
            O => \N__31102\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\
        );

    \I__4932\ : InMux
    port map (
            O => \N__31097\,
            I => \N__31093\
        );

    \I__4931\ : InMux
    port map (
            O => \N__31096\,
            I => \N__31090\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__31093\,
            I => \N__31087\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__31090\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_13\
        );

    \I__4928\ : Odrv4
    port map (
            O => \N__31087\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_13\
        );

    \I__4927\ : CascadeMux
    port map (
            O => \N__31082\,
            I => \N__31079\
        );

    \I__4926\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31076\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__31076\,
            I => \N__31073\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__31073\,
            I => \phase_controller_inst2.stoper_hc.counter_i_13\
        );

    \I__4923\ : InMux
    port map (
            O => \N__31070\,
            I => \N__31066\
        );

    \I__4922\ : InMux
    port map (
            O => \N__31069\,
            I => \N__31063\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__31066\,
            I => \N__31060\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__31063\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_14\
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__31060\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_14\
        );

    \I__4918\ : CascadeMux
    port map (
            O => \N__31055\,
            I => \N__31052\
        );

    \I__4917\ : InMux
    port map (
            O => \N__31052\,
            I => \N__31049\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__31049\,
            I => \phase_controller_inst2.stoper_hc.counter_i_14\
        );

    \I__4915\ : InMux
    port map (
            O => \N__31046\,
            I => \N__31042\
        );

    \I__4914\ : InMux
    port map (
            O => \N__31045\,
            I => \N__31039\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__31042\,
            I => \N__31036\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__31039\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_15\
        );

    \I__4911\ : Odrv4
    port map (
            O => \N__31036\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_15\
        );

    \I__4910\ : InMux
    port map (
            O => \N__31031\,
            I => \N__31028\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__31028\,
            I => \phase_controller_inst2.stoper_hc.counter_i_15\
        );

    \I__4908\ : InMux
    port map (
            O => \N__31025\,
            I => \N__31022\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__31022\,
            I => \N__31019\
        );

    \I__4906\ : Span4Mux_h
    port map (
            O => \N__31019\,
            I => \N__31016\
        );

    \I__4905\ : Odrv4
    port map (
            O => \N__31016\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt16\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__31013\,
            I => \N__31010\
        );

    \I__4903\ : InMux
    port map (
            O => \N__31010\,
            I => \N__31007\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__31007\,
            I => \N__31004\
        );

    \I__4901\ : Span4Mux_h
    port map (
            O => \N__31004\,
            I => \N__31001\
        );

    \I__4900\ : Odrv4
    port map (
            O => \N__31001\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16\
        );

    \I__4899\ : InMux
    port map (
            O => \N__30998\,
            I => \N__30995\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__30995\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18\
        );

    \I__4897\ : CascadeMux
    port map (
            O => \N__30992\,
            I => \N__30989\
        );

    \I__4896\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30986\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__30986\,
            I => \N__30983\
        );

    \I__4894\ : Span4Mux_h
    port map (
            O => \N__30983\,
            I => \N__30980\
        );

    \I__4893\ : Odrv4
    port map (
            O => \N__30980\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt18\
        );

    \I__4892\ : InMux
    port map (
            O => \N__30977\,
            I => \N__30974\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__30974\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt20\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__30971\,
            I => \N__30968\
        );

    \I__4889\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30965\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__30965\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20\
        );

    \I__4887\ : InMux
    port map (
            O => \N__30962\,
            I => \N__30959\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__30959\,
            I => \N__30956\
        );

    \I__4885\ : Odrv4
    port map (
            O => \N__30956\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__30953\,
            I => \N__30950\
        );

    \I__4883\ : InMux
    port map (
            O => \N__30950\,
            I => \N__30947\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__30947\,
            I => \N__30944\
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__30944\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt22\
        );

    \I__4880\ : InMux
    port map (
            O => \N__30941\,
            I => \N__30938\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__30938\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24\
        );

    \I__4878\ : CascadeMux
    port map (
            O => \N__30935\,
            I => \N__30932\
        );

    \I__4877\ : InMux
    port map (
            O => \N__30932\,
            I => \N__30929\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__30929\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt24\
        );

    \I__4875\ : InMux
    port map (
            O => \N__30926\,
            I => \N__30922\
        );

    \I__4874\ : InMux
    port map (
            O => \N__30925\,
            I => \N__30919\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__30922\,
            I => \N__30916\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__30919\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_5\
        );

    \I__4871\ : Odrv4
    port map (
            O => \N__30916\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_5\
        );

    \I__4870\ : InMux
    port map (
            O => \N__30911\,
            I => \N__30908\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__30908\,
            I => \phase_controller_inst2.stoper_hc.counter_i_5\
        );

    \I__4868\ : InMux
    port map (
            O => \N__30905\,
            I => \N__30901\
        );

    \I__4867\ : InMux
    port map (
            O => \N__30904\,
            I => \N__30898\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__30901\,
            I => \N__30895\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__30898\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_6\
        );

    \I__4864\ : Odrv4
    port map (
            O => \N__30895\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_6\
        );

    \I__4863\ : InMux
    port map (
            O => \N__30890\,
            I => \N__30887\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__30887\,
            I => \phase_controller_inst2.stoper_hc.counter_i_6\
        );

    \I__4861\ : InMux
    port map (
            O => \N__30884\,
            I => \N__30880\
        );

    \I__4860\ : InMux
    port map (
            O => \N__30883\,
            I => \N__30877\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__30880\,
            I => \N__30874\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__30877\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_7\
        );

    \I__4857\ : Odrv4
    port map (
            O => \N__30874\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_7\
        );

    \I__4856\ : InMux
    port map (
            O => \N__30869\,
            I => \N__30866\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__30866\,
            I => \phase_controller_inst2.stoper_hc.counter_i_7\
        );

    \I__4854\ : InMux
    port map (
            O => \N__30863\,
            I => \N__30860\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__30860\,
            I => \N__30856\
        );

    \I__4852\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30853\
        );

    \I__4851\ : Span4Mux_v
    port map (
            O => \N__30856\,
            I => \N__30850\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__30853\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_8\
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__30850\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_8\
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__30845\,
            I => \N__30842\
        );

    \I__4847\ : InMux
    port map (
            O => \N__30842\,
            I => \N__30839\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__30839\,
            I => \phase_controller_inst2.stoper_hc.counter_i_8\
        );

    \I__4845\ : InMux
    port map (
            O => \N__30836\,
            I => \N__30832\
        );

    \I__4844\ : InMux
    port map (
            O => \N__30835\,
            I => \N__30829\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__30832\,
            I => \N__30826\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__30829\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_9\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__30826\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_9\
        );

    \I__4840\ : InMux
    port map (
            O => \N__30821\,
            I => \N__30818\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__30818\,
            I => \phase_controller_inst2.stoper_hc.counter_i_9\
        );

    \I__4838\ : InMux
    port map (
            O => \N__30815\,
            I => \N__30812\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__30812\,
            I => \N__30808\
        );

    \I__4836\ : InMux
    port map (
            O => \N__30811\,
            I => \N__30805\
        );

    \I__4835\ : Span4Mux_v
    port map (
            O => \N__30808\,
            I => \N__30802\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__30805\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_10\
        );

    \I__4833\ : Odrv4
    port map (
            O => \N__30802\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_10\
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__30797\,
            I => \N__30794\
        );

    \I__4831\ : InMux
    port map (
            O => \N__30794\,
            I => \N__30791\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__30791\,
            I => \phase_controller_inst2.stoper_hc.counter_i_10\
        );

    \I__4829\ : InMux
    port map (
            O => \N__30788\,
            I => \N__30784\
        );

    \I__4828\ : InMux
    port map (
            O => \N__30787\,
            I => \N__30781\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__30784\,
            I => \N__30778\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__30781\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_11\
        );

    \I__4825\ : Odrv4
    port map (
            O => \N__30778\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_11\
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__30773\,
            I => \N__30770\
        );

    \I__4823\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30767\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__30767\,
            I => \N__30764\
        );

    \I__4821\ : Odrv4
    port map (
            O => \N__30764\,
            I => \phase_controller_inst2.stoper_hc.counter_i_11\
        );

    \I__4820\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30757\
        );

    \I__4819\ : InMux
    port map (
            O => \N__30760\,
            I => \N__30754\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__30757\,
            I => \N__30751\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__30754\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_12\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__30751\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_12\
        );

    \I__4815\ : CascadeMux
    port map (
            O => \N__30746\,
            I => \N__30743\
        );

    \I__4814\ : InMux
    port map (
            O => \N__30743\,
            I => \N__30740\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__30740\,
            I => \phase_controller_inst2.stoper_hc.counter_i_12\
        );

    \I__4812\ : InMux
    port map (
            O => \N__30737\,
            I => \N__30734\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__30734\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\
        );

    \I__4810\ : CascadeMux
    port map (
            O => \N__30731\,
            I => \N__30726\
        );

    \I__4809\ : InMux
    port map (
            O => \N__30730\,
            I => \N__30723\
        );

    \I__4808\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30717\
        );

    \I__4807\ : InMux
    port map (
            O => \N__30726\,
            I => \N__30717\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__30723\,
            I => \N__30714\
        );

    \I__4805\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30711\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__30717\,
            I => \N__30708\
        );

    \I__4803\ : Span12Mux_s11_v
    port map (
            O => \N__30714\,
            I => \N__30705\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__30711\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__4801\ : Odrv12
    port map (
            O => \N__30708\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__4800\ : Odrv12
    port map (
            O => \N__30705\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__4799\ : IoInMux
    port map (
            O => \N__30698\,
            I => \N__30695\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__30695\,
            I => \N__30692\
        );

    \I__4797\ : Span4Mux_s2_v
    port map (
            O => \N__30692\,
            I => \N__30689\
        );

    \I__4796\ : Odrv4
    port map (
            O => \N__30689\,
            I => s2_phy_c
        );

    \I__4795\ : InMux
    port map (
            O => \N__30686\,
            I => \N__30679\
        );

    \I__4794\ : CascadeMux
    port map (
            O => \N__30685\,
            I => \N__30676\
        );

    \I__4793\ : InMux
    port map (
            O => \N__30684\,
            I => \N__30672\
        );

    \I__4792\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30667\
        );

    \I__4791\ : InMux
    port map (
            O => \N__30682\,
            I => \N__30667\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__30679\,
            I => \N__30664\
        );

    \I__4789\ : InMux
    port map (
            O => \N__30676\,
            I => \N__30661\
        );

    \I__4788\ : InMux
    port map (
            O => \N__30675\,
            I => \N__30658\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__30672\,
            I => \N__30655\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__30667\,
            I => \N__30652\
        );

    \I__4785\ : Span12Mux_s6_v
    port map (
            O => \N__30664\,
            I => \N__30649\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__30661\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__30658\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__4782\ : Odrv12
    port map (
            O => \N__30655\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__4781\ : Odrv4
    port map (
            O => \N__30652\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__4780\ : Odrv12
    port map (
            O => \N__30649\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__4779\ : CascadeMux
    port map (
            O => \N__30638\,
            I => \N__30634\
        );

    \I__4778\ : InMux
    port map (
            O => \N__30637\,
            I => \N__30631\
        );

    \I__4777\ : InMux
    port map (
            O => \N__30634\,
            I => \N__30628\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__30631\,
            I => \phase_controller_inst2.stoper_hc.counter\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__30628\,
            I => \phase_controller_inst2.stoper_hc.counter\
        );

    \I__4774\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30620\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__30620\,
            I => \N__30616\
        );

    \I__4772\ : InMux
    port map (
            O => \N__30619\,
            I => \N__30613\
        );

    \I__4771\ : Span4Mux_v
    port map (
            O => \N__30616\,
            I => \N__30610\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__30613\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_0\
        );

    \I__4769\ : Odrv4
    port map (
            O => \N__30610\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_0\
        );

    \I__4768\ : InMux
    port map (
            O => \N__30605\,
            I => \N__30602\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__30602\,
            I => \phase_controller_inst2.stoper_hc.counter_i_0\
        );

    \I__4766\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30595\
        );

    \I__4765\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30592\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__30595\,
            I => \N__30589\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__30592\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_1\
        );

    \I__4762\ : Odrv4
    port map (
            O => \N__30589\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_1\
        );

    \I__4761\ : CascadeMux
    port map (
            O => \N__30584\,
            I => \N__30581\
        );

    \I__4760\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30578\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__30578\,
            I => \phase_controller_inst2.stoper_hc.counter_i_1\
        );

    \I__4758\ : InMux
    port map (
            O => \N__30575\,
            I => \N__30572\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__30572\,
            I => \N__30568\
        );

    \I__4756\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30565\
        );

    \I__4755\ : Span4Mux_v
    port map (
            O => \N__30568\,
            I => \N__30562\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__30565\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_2\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__30562\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_2\
        );

    \I__4752\ : CascadeMux
    port map (
            O => \N__30557\,
            I => \N__30554\
        );

    \I__4751\ : InMux
    port map (
            O => \N__30554\,
            I => \N__30551\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__30551\,
            I => \phase_controller_inst2.stoper_hc.counter_i_2\
        );

    \I__4749\ : InMux
    port map (
            O => \N__30548\,
            I => \N__30544\
        );

    \I__4748\ : InMux
    port map (
            O => \N__30547\,
            I => \N__30541\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__30544\,
            I => \N__30538\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__30541\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_3\
        );

    \I__4745\ : Odrv4
    port map (
            O => \N__30538\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_3\
        );

    \I__4744\ : InMux
    port map (
            O => \N__30533\,
            I => \N__30530\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__30530\,
            I => \phase_controller_inst2.stoper_hc.counter_i_3\
        );

    \I__4742\ : InMux
    port map (
            O => \N__30527\,
            I => \N__30523\
        );

    \I__4741\ : InMux
    port map (
            O => \N__30526\,
            I => \N__30520\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__30523\,
            I => \N__30517\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__30520\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_4\
        );

    \I__4738\ : Odrv4
    port map (
            O => \N__30517\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_4\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__30512\,
            I => \N__30509\
        );

    \I__4736\ : InMux
    port map (
            O => \N__30509\,
            I => \N__30506\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__30506\,
            I => \phase_controller_inst2.stoper_hc.counter_i_4\
        );

    \I__4734\ : InMux
    port map (
            O => \N__30503\,
            I => \N__30500\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__30500\,
            I => \N__30496\
        );

    \I__4732\ : InMux
    port map (
            O => \N__30499\,
            I => \N__30493\
        );

    \I__4731\ : Odrv4
    port map (
            O => \N__30496\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__30493\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21\
        );

    \I__4729\ : InMux
    port map (
            O => \N__30488\,
            I => \N__30484\
        );

    \I__4728\ : InMux
    port map (
            O => \N__30487\,
            I => \N__30481\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__30484\,
            I => \N__30477\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__30481\,
            I => \N__30474\
        );

    \I__4725\ : InMux
    port map (
            O => \N__30480\,
            I => \N__30471\
        );

    \I__4724\ : Span4Mux_v
    port map (
            O => \N__30477\,
            I => \N__30466\
        );

    \I__4723\ : Span4Mux_v
    port map (
            O => \N__30474\,
            I => \N__30466\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__30471\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_21\
        );

    \I__4721\ : Odrv4
    port map (
            O => \N__30466\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_21\
        );

    \I__4720\ : CascadeMux
    port map (
            O => \N__30461\,
            I => \N__30458\
        );

    \I__4719\ : InMux
    port map (
            O => \N__30458\,
            I => \N__30454\
        );

    \I__4718\ : InMux
    port map (
            O => \N__30457\,
            I => \N__30451\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__30454\,
            I => \N__30448\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__30451\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20\
        );

    \I__4715\ : Odrv4
    port map (
            O => \N__30448\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20\
        );

    \I__4714\ : CascadeMux
    port map (
            O => \N__30443\,
            I => \N__30439\
        );

    \I__4713\ : InMux
    port map (
            O => \N__30442\,
            I => \N__30436\
        );

    \I__4712\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30433\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__30436\,
            I => \N__30427\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__30433\,
            I => \N__30427\
        );

    \I__4709\ : InMux
    port map (
            O => \N__30432\,
            I => \N__30424\
        );

    \I__4708\ : Span4Mux_v
    port map (
            O => \N__30427\,
            I => \N__30421\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__30424\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_20\
        );

    \I__4706\ : Odrv4
    port map (
            O => \N__30421\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_20\
        );

    \I__4705\ : InMux
    port map (
            O => \N__30416\,
            I => \N__30413\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__30413\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt20\
        );

    \I__4703\ : InMux
    port map (
            O => \N__30410\,
            I => \N__30407\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__30407\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__4701\ : CascadeMux
    port map (
            O => \N__30404\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\
        );

    \I__4700\ : InMux
    port map (
            O => \N__30401\,
            I => \N__30398\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__30398\,
            I => \N__30395\
        );

    \I__4698\ : Span4Mux_h
    port map (
            O => \N__30395\,
            I => \N__30392\
        );

    \I__4697\ : Span4Mux_v
    port map (
            O => \N__30392\,
            I => \N__30389\
        );

    \I__4696\ : Odrv4
    port map (
            O => \N__30389\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19\
        );

    \I__4695\ : InMux
    port map (
            O => \N__30386\,
            I => \N__30382\
        );

    \I__4694\ : InMux
    port map (
            O => \N__30385\,
            I => \N__30379\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__30382\,
            I => \N__30374\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__30379\,
            I => \N__30374\
        );

    \I__4691\ : Odrv4
    port map (
            O => \N__30374\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_22\
        );

    \I__4690\ : InMux
    port map (
            O => \N__30371\,
            I => \N__30368\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__30368\,
            I => \N__30364\
        );

    \I__4688\ : InMux
    port map (
            O => \N__30367\,
            I => \N__30360\
        );

    \I__4687\ : Span4Mux_h
    port map (
            O => \N__30364\,
            I => \N__30357\
        );

    \I__4686\ : InMux
    port map (
            O => \N__30363\,
            I => \N__30354\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__30360\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_23\
        );

    \I__4684\ : Odrv4
    port map (
            O => \N__30357\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_23\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__30354\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_23\
        );

    \I__4682\ : CascadeMux
    port map (
            O => \N__30347\,
            I => \N__30344\
        );

    \I__4681\ : InMux
    port map (
            O => \N__30344\,
            I => \N__30340\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__30343\,
            I => \N__30336\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__30340\,
            I => \N__30333\
        );

    \I__4678\ : InMux
    port map (
            O => \N__30339\,
            I => \N__30330\
        );

    \I__4677\ : InMux
    port map (
            O => \N__30336\,
            I => \N__30327\
        );

    \I__4676\ : Span4Mux_h
    port map (
            O => \N__30333\,
            I => \N__30324\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__30330\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_22\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__30327\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_22\
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__30324\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_22\
        );

    \I__4672\ : InMux
    port map (
            O => \N__30317\,
            I => \N__30313\
        );

    \I__4671\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30310\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__30313\,
            I => \N__30305\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__30310\,
            I => \N__30305\
        );

    \I__4668\ : Odrv4
    port map (
            O => \N__30305\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_23\
        );

    \I__4667\ : CascadeMux
    port map (
            O => \N__30302\,
            I => \N__30299\
        );

    \I__4666\ : InMux
    port map (
            O => \N__30299\,
            I => \N__30296\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__30296\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt22\
        );

    \I__4664\ : InMux
    port map (
            O => \N__30293\,
            I => \N__30290\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__30290\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\
        );

    \I__4662\ : CascadeMux
    port map (
            O => \N__30287\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_\
        );

    \I__4661\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30281\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__30281\,
            I => \N__30278\
        );

    \I__4659\ : Span12Mux_v
    port map (
            O => \N__30278\,
            I => \N__30275\
        );

    \I__4658\ : Odrv12
    port map (
            O => \N__30275\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\
        );

    \I__4657\ : InMux
    port map (
            O => \N__30272\,
            I => \N__30269\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__30269\,
            I => \N__30266\
        );

    \I__4655\ : Span4Mux_h
    port map (
            O => \N__30266\,
            I => \N__30263\
        );

    \I__4654\ : Sp12to4
    port map (
            O => \N__30263\,
            I => \N__30260\
        );

    \I__4653\ : Span12Mux_v
    port map (
            O => \N__30260\,
            I => \N__30257\
        );

    \I__4652\ : Odrv12
    port map (
            O => \N__30257\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_15\
        );

    \I__4651\ : InMux
    port map (
            O => \N__30254\,
            I => \N__30251\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__30251\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\
        );

    \I__4649\ : CascadeMux
    port map (
            O => \N__30248\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\
        );

    \I__4648\ : InMux
    port map (
            O => \N__30245\,
            I => \N__30242\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__30242\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28\
        );

    \I__4646\ : InMux
    port map (
            O => \N__30239\,
            I => \N__30235\
        );

    \I__4645\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30232\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__30235\,
            I => \N__30229\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__30232\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_20
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__30229\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_20
        );

    \I__4641\ : InMux
    port map (
            O => \N__30224\,
            I => \N__30220\
        );

    \I__4640\ : InMux
    port map (
            O => \N__30223\,
            I => \N__30217\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__30220\,
            I => \N__30214\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__30217\,
            I => \N__30211\
        );

    \I__4637\ : Odrv4
    port map (
            O => \N__30214\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_21
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__30211\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_21
        );

    \I__4635\ : InMux
    port map (
            O => \N__30206\,
            I => \N__30202\
        );

    \I__4634\ : InMux
    port map (
            O => \N__30205\,
            I => \N__30199\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__30202\,
            I => \N__30196\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__30199\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_22
        );

    \I__4631\ : Odrv4
    port map (
            O => \N__30196\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_22
        );

    \I__4630\ : InMux
    port map (
            O => \N__30191\,
            I => \N__30188\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__30188\,
            I => \N__30185\
        );

    \I__4628\ : Span4Mux_v
    port map (
            O => \N__30185\,
            I => \N__30181\
        );

    \I__4627\ : InMux
    port map (
            O => \N__30184\,
            I => \N__30178\
        );

    \I__4626\ : Span4Mux_v
    port map (
            O => \N__30181\,
            I => \N__30173\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__30178\,
            I => \N__30173\
        );

    \I__4624\ : Odrv4
    port map (
            O => \N__30173\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_23
        );

    \I__4623\ : CascadeMux
    port map (
            O => \N__30170\,
            I => \N__30167\
        );

    \I__4622\ : InMux
    port map (
            O => \N__30167\,
            I => \N__30164\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__30164\,
            I => \N__30161\
        );

    \I__4620\ : Odrv4
    port map (
            O => \N__30161\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20\
        );

    \I__4619\ : InMux
    port map (
            O => \N__30158\,
            I => \N__30155\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__30155\,
            I => \N__30152\
        );

    \I__4617\ : Span4Mux_v
    port map (
            O => \N__30152\,
            I => \N__30149\
        );

    \I__4616\ : Odrv4
    port map (
            O => \N__30149\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\
        );

    \I__4615\ : CascadeMux
    port map (
            O => \N__30146\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\
        );

    \I__4614\ : InMux
    port map (
            O => \N__30143\,
            I => \N__30140\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__30140\,
            I => \N__30137\
        );

    \I__4612\ : Odrv12
    port map (
            O => \N__30137\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\
        );

    \I__4611\ : InMux
    port map (
            O => \N__30134\,
            I => \N__30131\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__30131\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26\
        );

    \I__4609\ : InMux
    port map (
            O => \N__30128\,
            I => \N__30125\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__30125\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__4607\ : CascadeMux
    port map (
            O => \N__30122\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\
        );

    \I__4606\ : InMux
    port map (
            O => \N__30119\,
            I => \N__30116\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__30116\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18\
        );

    \I__4604\ : InMux
    port map (
            O => \N__30113\,
            I => \N__30109\
        );

    \I__4603\ : InMux
    port map (
            O => \N__30112\,
            I => \N__30106\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__30109\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__30106\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__4600\ : InMux
    port map (
            O => \N__30101\,
            I => \N__30098\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__30098\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__4598\ : CascadeMux
    port map (
            O => \N__30095\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\
        );

    \I__4597\ : InMux
    port map (
            O => \N__30092\,
            I => \N__30089\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__30089\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27\
        );

    \I__4595\ : InMux
    port map (
            O => \N__30086\,
            I => \N__30083\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__30083\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__4593\ : CascadeMux
    port map (
            O => \N__30080\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\
        );

    \I__4592\ : InMux
    port map (
            O => \N__30077\,
            I => \N__30074\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__30074\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25\
        );

    \I__4590\ : InMux
    port map (
            O => \N__30071\,
            I => \N__30068\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__30068\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__4588\ : CascadeMux
    port map (
            O => \N__30065\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\
        );

    \I__4587\ : InMux
    port map (
            O => \N__30062\,
            I => \N__30059\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__30059\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16\
        );

    \I__4585\ : InMux
    port map (
            O => \N__30056\,
            I => \N__30052\
        );

    \I__4584\ : InMux
    port map (
            O => \N__30055\,
            I => \N__30049\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__30052\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__30049\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4581\ : InMux
    port map (
            O => \N__30044\,
            I => \N__30041\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__30041\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12\
        );

    \I__4579\ : InMux
    port map (
            O => \N__30038\,
            I => \N__30035\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__30035\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__4577\ : CascadeMux
    port map (
            O => \N__30032\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\
        );

    \I__4576\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30026\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__30026\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10\
        );

    \I__4574\ : InMux
    port map (
            O => \N__30023\,
            I => \N__30020\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__30020\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__30017\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17_cascade_\
        );

    \I__4571\ : CascadeMux
    port map (
            O => \N__30014\,
            I => \N__30011\
        );

    \I__4570\ : InMux
    port map (
            O => \N__30011\,
            I => \N__30008\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__30008\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17\
        );

    \I__4568\ : InMux
    port map (
            O => \N__30005\,
            I => \N__30001\
        );

    \I__4567\ : InMux
    port map (
            O => \N__30004\,
            I => \N__29998\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__30001\,
            I => \N__29995\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__29998\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__4564\ : Odrv12
    port map (
            O => \N__29995\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__4563\ : InMux
    port map (
            O => \N__29990\,
            I => \N__29987\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__29987\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30\
        );

    \I__4561\ : InMux
    port map (
            O => \N__29984\,
            I => \N__29981\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__29981\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__4559\ : CascadeMux
    port map (
            O => \N__29978\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\
        );

    \I__4558\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29972\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__29972\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__29969\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4_cascade_\
        );

    \I__4555\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29963\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__29963\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4\
        );

    \I__4553\ : InMux
    port map (
            O => \N__29960\,
            I => \N__29956\
        );

    \I__4552\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29953\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__29956\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__29953\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__4549\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29945\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__29945\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11\
        );

    \I__4547\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29939\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__29939\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__4545\ : CascadeMux
    port map (
            O => \N__29936\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\
        );

    \I__4544\ : CascadeMux
    port map (
            O => \N__29933\,
            I => \N__29930\
        );

    \I__4543\ : InMux
    port map (
            O => \N__29930\,
            I => \N__29927\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__29927\,
            I => \N__29924\
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__29924\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20\
        );

    \I__4540\ : InMux
    port map (
            O => \N__29921\,
            I => \N__29917\
        );

    \I__4539\ : InMux
    port map (
            O => \N__29920\,
            I => \N__29914\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__29917\,
            I => \N__29911\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__29914\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__4536\ : Odrv4
    port map (
            O => \N__29911\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__4535\ : InMux
    port map (
            O => \N__29906\,
            I => \N__29903\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__29903\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24\
        );

    \I__4533\ : InMux
    port map (
            O => \N__29900\,
            I => \N__29897\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__29897\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__4531\ : CascadeMux
    port map (
            O => \N__29894\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5_cascade_\
        );

    \I__4530\ : InMux
    port map (
            O => \N__29891\,
            I => \N__29888\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__29888\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5\
        );

    \I__4528\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29882\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__29882\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__4526\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29875\
        );

    \I__4525\ : InMux
    port map (
            O => \N__29878\,
            I => \N__29872\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__29875\,
            I => \N__29869\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__29872\,
            I => \N__29866\
        );

    \I__4522\ : Span12Mux_v
    port map (
            O => \N__29869\,
            I => \N__29863\
        );

    \I__4521\ : Span12Mux_v
    port map (
            O => \N__29866\,
            I => \N__29860\
        );

    \I__4520\ : Span12Mux_h
    port map (
            O => \N__29863\,
            I => \N__29857\
        );

    \I__4519\ : Span12Mux_h
    port map (
            O => \N__29860\,
            I => \N__29854\
        );

    \I__4518\ : Span12Mux_h
    port map (
            O => \N__29857\,
            I => \N__29851\
        );

    \I__4517\ : Odrv12
    port map (
            O => \N__29854\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__4516\ : Odrv12
    port map (
            O => \N__29851\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__4515\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29843\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__29843\,
            I => \N__29840\
        );

    \I__4513\ : Span4Mux_h
    port map (
            O => \N__29840\,
            I => \N__29837\
        );

    \I__4512\ : Sp12to4
    port map (
            O => \N__29837\,
            I => \N__29834\
        );

    \I__4511\ : Span12Mux_v
    port map (
            O => \N__29834\,
            I => \N__29831\
        );

    \I__4510\ : Odrv12
    port map (
            O => \N__29831\,
            I => \pwm_generator_inst.un3_threshold_iZ0\
        );

    \I__4509\ : InMux
    port map (
            O => \N__29828\,
            I => \N__29825\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__29825\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\
        );

    \I__4507\ : CascadeMux
    port map (
            O => \N__29822\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\
        );

    \I__4506\ : CascadeMux
    port map (
            O => \N__29819\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\
        );

    \I__4505\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29813\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__29813\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4503\ : CascadeMux
    port map (
            O => \N__29810\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6_cascade_\
        );

    \I__4502\ : InMux
    port map (
            O => \N__29807\,
            I => \N__29804\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__29804\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6\
        );

    \I__4500\ : InMux
    port map (
            O => \N__29801\,
            I => \N__29798\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__29798\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__4498\ : CascadeMux
    port map (
            O => \N__29795\,
            I => \elapsed_time_ns_1_RNILK91B_0_9_cascade_\
        );

    \I__4497\ : InMux
    port map (
            O => \N__29792\,
            I => \N__29789\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__29789\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9\
        );

    \I__4495\ : InMux
    port map (
            O => \N__29786\,
            I => \N__29782\
        );

    \I__4494\ : InMux
    port map (
            O => \N__29785\,
            I => \N__29779\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__29782\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__29779\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__4491\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29764\
        );

    \I__4490\ : InMux
    port map (
            O => \N__29773\,
            I => \N__29764\
        );

    \I__4489\ : InMux
    port map (
            O => \N__29772\,
            I => \N__29764\
        );

    \I__4488\ : InMux
    port map (
            O => \N__29771\,
            I => \N__29761\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__29764\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__29761\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__4485\ : InMux
    port map (
            O => \N__29756\,
            I => \N__29753\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__29753\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa\
        );

    \I__4483\ : InMux
    port map (
            O => \N__29750\,
            I => \N__29747\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__29747\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__29744\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\
        );

    \I__4480\ : InMux
    port map (
            O => \N__29741\,
            I => \N__29738\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__29738\,
            I => \N__29735\
        );

    \I__4478\ : Odrv4
    port map (
            O => \N__29735\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13\
        );

    \I__4477\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29729\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__29729\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__4475\ : CascadeMux
    port map (
            O => \N__29726\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8_cascade_\
        );

    \I__4474\ : InMux
    port map (
            O => \N__29723\,
            I => \N__29720\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__29720\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8\
        );

    \I__4472\ : InMux
    port map (
            O => \N__29717\,
            I => \N__29710\
        );

    \I__4471\ : InMux
    port map (
            O => \N__29716\,
            I => \N__29710\
        );

    \I__4470\ : InMux
    port map (
            O => \N__29715\,
            I => \N__29707\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__29710\,
            I => \N__29704\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__29707\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_17\
        );

    \I__4467\ : Odrv12
    port map (
            O => \N__29704\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_17\
        );

    \I__4466\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29693\
        );

    \I__4465\ : InMux
    port map (
            O => \N__29698\,
            I => \N__29693\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__29693\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_16\
        );

    \I__4463\ : CascadeMux
    port map (
            O => \N__29690\,
            I => \N__29686\
        );

    \I__4462\ : CascadeMux
    port map (
            O => \N__29689\,
            I => \N__29683\
        );

    \I__4461\ : InMux
    port map (
            O => \N__29686\,
            I => \N__29677\
        );

    \I__4460\ : InMux
    port map (
            O => \N__29683\,
            I => \N__29677\
        );

    \I__4459\ : InMux
    port map (
            O => \N__29682\,
            I => \N__29674\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__29677\,
            I => \N__29671\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__29674\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_16\
        );

    \I__4456\ : Odrv12
    port map (
            O => \N__29671\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_16\
        );

    \I__4455\ : InMux
    port map (
            O => \N__29666\,
            I => \N__29662\
        );

    \I__4454\ : InMux
    port map (
            O => \N__29665\,
            I => \N__29659\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__29662\,
            I => \N__29656\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__29659\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18\
        );

    \I__4451\ : Odrv4
    port map (
            O => \N__29656\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18\
        );

    \I__4450\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29639\
        );

    \I__4449\ : InMux
    port map (
            O => \N__29650\,
            I => \N__29639\
        );

    \I__4448\ : InMux
    port map (
            O => \N__29649\,
            I => \N__29639\
        );

    \I__4447\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29639\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__29639\,
            I => \N__29636\
        );

    \I__4445\ : Span4Mux_h
    port map (
            O => \N__29636\,
            I => \N__29633\
        );

    \I__4444\ : Odrv4
    port map (
            O => \N__29633\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28\
        );

    \I__4443\ : InMux
    port map (
            O => \N__29630\,
            I => \N__29624\
        );

    \I__4442\ : InMux
    port map (
            O => \N__29629\,
            I => \N__29624\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__29624\,
            I => \N__29621\
        );

    \I__4440\ : Odrv12
    port map (
            O => \N__29621\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_26\
        );

    \I__4439\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29615\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__29615\,
            I => \N__29610\
        );

    \I__4437\ : InMux
    port map (
            O => \N__29614\,
            I => \N__29607\
        );

    \I__4436\ : InMux
    port map (
            O => \N__29613\,
            I => \N__29604\
        );

    \I__4435\ : Span12Mux_h
    port map (
            O => \N__29610\,
            I => \N__29597\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__29607\,
            I => \N__29597\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__29604\,
            I => \N__29597\
        );

    \I__4432\ : Odrv12
    port map (
            O => \N__29597\,
            I => il_min_comp1_c
        );

    \I__4431\ : InMux
    port map (
            O => \N__29594\,
            I => \N__29587\
        );

    \I__4430\ : InMux
    port map (
            O => \N__29593\,
            I => \N__29587\
        );

    \I__4429\ : InMux
    port map (
            O => \N__29592\,
            I => \N__29584\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__29587\,
            I => \N__29579\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__29584\,
            I => \N__29579\
        );

    \I__4426\ : Span4Mux_h
    port map (
            O => \N__29579\,
            I => \N__29576\
        );

    \I__4425\ : Span4Mux_v
    port map (
            O => \N__29576\,
            I => \N__29573\
        );

    \I__4424\ : Span4Mux_v
    port map (
            O => \N__29573\,
            I => \N__29570\
        );

    \I__4423\ : Odrv4
    port map (
            O => \N__29570\,
            I => il_max_comp1_c
        );

    \I__4422\ : InMux
    port map (
            O => \N__29567\,
            I => \N__29560\
        );

    \I__4421\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29560\
        );

    \I__4420\ : InMux
    port map (
            O => \N__29565\,
            I => \N__29557\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__29560\,
            I => \N__29554\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__29557\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_25\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__29554\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_25\
        );

    \I__4416\ : InMux
    port map (
            O => \N__29549\,
            I => \N__29542\
        );

    \I__4415\ : InMux
    port map (
            O => \N__29548\,
            I => \N__29542\
        );

    \I__4414\ : InMux
    port map (
            O => \N__29547\,
            I => \N__29539\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__29542\,
            I => \N__29536\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__29539\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_24\
        );

    \I__4411\ : Odrv4
    port map (
            O => \N__29536\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_24\
        );

    \I__4410\ : InMux
    port map (
            O => \N__29531\,
            I => \N__29524\
        );

    \I__4409\ : InMux
    port map (
            O => \N__29530\,
            I => \N__29524\
        );

    \I__4408\ : InMux
    port map (
            O => \N__29529\,
            I => \N__29521\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__29524\,
            I => \N__29518\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__29521\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_27\
        );

    \I__4405\ : Odrv4
    port map (
            O => \N__29518\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_27\
        );

    \I__4404\ : InMux
    port map (
            O => \N__29513\,
            I => \N__29506\
        );

    \I__4403\ : InMux
    port map (
            O => \N__29512\,
            I => \N__29506\
        );

    \I__4402\ : InMux
    port map (
            O => \N__29511\,
            I => \N__29503\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__29506\,
            I => \N__29500\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__29503\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_26\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__29500\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_26\
        );

    \I__4398\ : CascadeMux
    port map (
            O => \N__29495\,
            I => \N__29492\
        );

    \I__4397\ : InMux
    port map (
            O => \N__29492\,
            I => \N__29487\
        );

    \I__4396\ : InMux
    port map (
            O => \N__29491\,
            I => \N__29484\
        );

    \I__4395\ : InMux
    port map (
            O => \N__29490\,
            I => \N__29481\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__29487\,
            I => \N__29476\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__29484\,
            I => \N__29476\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__29481\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_18\
        );

    \I__4391\ : Odrv12
    port map (
            O => \N__29476\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_18\
        );

    \I__4390\ : CascadeMux
    port map (
            O => \N__29471\,
            I => \N__29468\
        );

    \I__4389\ : InMux
    port map (
            O => \N__29468\,
            I => \N__29464\
        );

    \I__4388\ : InMux
    port map (
            O => \N__29467\,
            I => \N__29460\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__29464\,
            I => \N__29457\
        );

    \I__4386\ : InMux
    port map (
            O => \N__29463\,
            I => \N__29454\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__29460\,
            I => \N__29451\
        );

    \I__4384\ : Span4Mux_v
    port map (
            O => \N__29457\,
            I => \N__29448\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__29454\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_19\
        );

    \I__4382\ : Odrv4
    port map (
            O => \N__29451\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_19\
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__29448\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_19\
        );

    \I__4380\ : InMux
    port map (
            O => \N__29441\,
            I => \N__29434\
        );

    \I__4379\ : InMux
    port map (
            O => \N__29440\,
            I => \N__29434\
        );

    \I__4378\ : InMux
    port map (
            O => \N__29439\,
            I => \N__29431\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__29434\,
            I => \N__29428\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__29431\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_22\
        );

    \I__4375\ : Odrv12
    port map (
            O => \N__29428\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_22\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__29423\,
            I => \N__29419\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__29422\,
            I => \N__29416\
        );

    \I__4372\ : InMux
    port map (
            O => \N__29419\,
            I => \N__29410\
        );

    \I__4371\ : InMux
    port map (
            O => \N__29416\,
            I => \N__29410\
        );

    \I__4370\ : InMux
    port map (
            O => \N__29415\,
            I => \N__29407\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__29410\,
            I => \N__29404\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__29407\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_23\
        );

    \I__4367\ : Odrv12
    port map (
            O => \N__29404\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_23\
        );

    \I__4366\ : InMux
    port map (
            O => \N__29399\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_28\
        );

    \I__4365\ : InMux
    port map (
            O => \N__29396\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_29\
        );

    \I__4364\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29369\
        );

    \I__4363\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29369\
        );

    \I__4362\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29369\
        );

    \I__4361\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29369\
        );

    \I__4360\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29360\
        );

    \I__4359\ : InMux
    port map (
            O => \N__29388\,
            I => \N__29360\
        );

    \I__4358\ : InMux
    port map (
            O => \N__29387\,
            I => \N__29360\
        );

    \I__4357\ : InMux
    port map (
            O => \N__29386\,
            I => \N__29360\
        );

    \I__4356\ : InMux
    port map (
            O => \N__29385\,
            I => \N__29337\
        );

    \I__4355\ : InMux
    port map (
            O => \N__29384\,
            I => \N__29337\
        );

    \I__4354\ : InMux
    port map (
            O => \N__29383\,
            I => \N__29337\
        );

    \I__4353\ : InMux
    port map (
            O => \N__29382\,
            I => \N__29326\
        );

    \I__4352\ : InMux
    port map (
            O => \N__29381\,
            I => \N__29326\
        );

    \I__4351\ : InMux
    port map (
            O => \N__29380\,
            I => \N__29326\
        );

    \I__4350\ : InMux
    port map (
            O => \N__29379\,
            I => \N__29326\
        );

    \I__4349\ : InMux
    port map (
            O => \N__29378\,
            I => \N__29326\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__29369\,
            I => \N__29323\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__29360\,
            I => \N__29320\
        );

    \I__4346\ : InMux
    port map (
            O => \N__29359\,
            I => \N__29311\
        );

    \I__4345\ : InMux
    port map (
            O => \N__29358\,
            I => \N__29311\
        );

    \I__4344\ : InMux
    port map (
            O => \N__29357\,
            I => \N__29311\
        );

    \I__4343\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29311\
        );

    \I__4342\ : InMux
    port map (
            O => \N__29355\,
            I => \N__29302\
        );

    \I__4341\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29302\
        );

    \I__4340\ : InMux
    port map (
            O => \N__29353\,
            I => \N__29302\
        );

    \I__4339\ : InMux
    port map (
            O => \N__29352\,
            I => \N__29302\
        );

    \I__4338\ : InMux
    port map (
            O => \N__29351\,
            I => \N__29293\
        );

    \I__4337\ : InMux
    port map (
            O => \N__29350\,
            I => \N__29293\
        );

    \I__4336\ : InMux
    port map (
            O => \N__29349\,
            I => \N__29293\
        );

    \I__4335\ : InMux
    port map (
            O => \N__29348\,
            I => \N__29293\
        );

    \I__4334\ : InMux
    port map (
            O => \N__29347\,
            I => \N__29284\
        );

    \I__4333\ : InMux
    port map (
            O => \N__29346\,
            I => \N__29284\
        );

    \I__4332\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29284\
        );

    \I__4331\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29284\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__29337\,
            I => \N__29279\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__29326\,
            I => \N__29279\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__29323\,
            I => \phase_controller_inst2.stoper_hc.start_latched_i_0\
        );

    \I__4327\ : Odrv4
    port map (
            O => \N__29320\,
            I => \phase_controller_inst2.stoper_hc.start_latched_i_0\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__29311\,
            I => \phase_controller_inst2.stoper_hc.start_latched_i_0\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__29302\,
            I => \phase_controller_inst2.stoper_hc.start_latched_i_0\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__29293\,
            I => \phase_controller_inst2.stoper_hc.start_latched_i_0\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__29284\,
            I => \phase_controller_inst2.stoper_hc.start_latched_i_0\
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__29279\,
            I => \phase_controller_inst2.stoper_hc.start_latched_i_0\
        );

    \I__4321\ : InMux
    port map (
            O => \N__29264\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_30\
        );

    \I__4320\ : CEMux
    port map (
            O => \N__29261\,
            I => \N__29257\
        );

    \I__4319\ : CEMux
    port map (
            O => \N__29260\,
            I => \N__29253\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__29257\,
            I => \N__29250\
        );

    \I__4317\ : CEMux
    port map (
            O => \N__29256\,
            I => \N__29246\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__29253\,
            I => \N__29241\
        );

    \I__4315\ : Span4Mux_v
    port map (
            O => \N__29250\,
            I => \N__29241\
        );

    \I__4314\ : CEMux
    port map (
            O => \N__29249\,
            I => \N__29238\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__29246\,
            I => \N__29233\
        );

    \I__4312\ : Span4Mux_s1_v
    port map (
            O => \N__29241\,
            I => \N__29233\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__29238\,
            I => \N__29230\
        );

    \I__4310\ : Odrv4
    port map (
            O => \N__29233\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__29230\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__4308\ : InMux
    port map (
            O => \N__29225\,
            I => \N__29220\
        );

    \I__4307\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29215\
        );

    \I__4306\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29215\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__29220\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_28\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__29215\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_28\
        );

    \I__4303\ : InMux
    port map (
            O => \N__29210\,
            I => \N__29205\
        );

    \I__4302\ : InMux
    port map (
            O => \N__29209\,
            I => \N__29200\
        );

    \I__4301\ : InMux
    port map (
            O => \N__29208\,
            I => \N__29200\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__29205\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_29\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__29200\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_29\
        );

    \I__4298\ : InMux
    port map (
            O => \N__29195\,
            I => \N__29190\
        );

    \I__4297\ : InMux
    port map (
            O => \N__29194\,
            I => \N__29185\
        );

    \I__4296\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29185\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__29190\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_30\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__29185\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_30\
        );

    \I__4293\ : InMux
    port map (
            O => \N__29180\,
            I => \N__29175\
        );

    \I__4292\ : InMux
    port map (
            O => \N__29179\,
            I => \N__29172\
        );

    \I__4291\ : InMux
    port map (
            O => \N__29178\,
            I => \N__29169\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__29175\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_31\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__29172\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_31\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__29169\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_31\
        );

    \I__4287\ : InMux
    port map (
            O => \N__29162\,
            I => \N__29155\
        );

    \I__4286\ : InMux
    port map (
            O => \N__29161\,
            I => \N__29155\
        );

    \I__4285\ : InMux
    port map (
            O => \N__29160\,
            I => \N__29152\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__29155\,
            I => \N__29149\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__29152\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_21\
        );

    \I__4282\ : Odrv4
    port map (
            O => \N__29149\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_21\
        );

    \I__4281\ : CascadeMux
    port map (
            O => \N__29144\,
            I => \N__29140\
        );

    \I__4280\ : CascadeMux
    port map (
            O => \N__29143\,
            I => \N__29137\
        );

    \I__4279\ : InMux
    port map (
            O => \N__29140\,
            I => \N__29131\
        );

    \I__4278\ : InMux
    port map (
            O => \N__29137\,
            I => \N__29131\
        );

    \I__4277\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29128\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__29131\,
            I => \N__29125\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__29128\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_20\
        );

    \I__4274\ : Odrv4
    port map (
            O => \N__29125\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_20\
        );

    \I__4273\ : InMux
    port map (
            O => \N__29120\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_19\
        );

    \I__4272\ : InMux
    port map (
            O => \N__29117\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_20\
        );

    \I__4271\ : InMux
    port map (
            O => \N__29114\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_21\
        );

    \I__4270\ : InMux
    port map (
            O => \N__29111\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_22\
        );

    \I__4269\ : InMux
    port map (
            O => \N__29108\,
            I => \bfn_10_5_0_\
        );

    \I__4268\ : InMux
    port map (
            O => \N__29105\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_24\
        );

    \I__4267\ : InMux
    port map (
            O => \N__29102\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_25\
        );

    \I__4266\ : InMux
    port map (
            O => \N__29099\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_26\
        );

    \I__4265\ : InMux
    port map (
            O => \N__29096\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_27\
        );

    \I__4264\ : InMux
    port map (
            O => \N__29093\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_10\
        );

    \I__4263\ : InMux
    port map (
            O => \N__29090\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_11\
        );

    \I__4262\ : InMux
    port map (
            O => \N__29087\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_12\
        );

    \I__4261\ : InMux
    port map (
            O => \N__29084\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_13\
        );

    \I__4260\ : InMux
    port map (
            O => \N__29081\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_14\
        );

    \I__4259\ : InMux
    port map (
            O => \N__29078\,
            I => \bfn_10_4_0_\
        );

    \I__4258\ : InMux
    port map (
            O => \N__29075\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_16\
        );

    \I__4257\ : InMux
    port map (
            O => \N__29072\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_17\
        );

    \I__4256\ : InMux
    port map (
            O => \N__29069\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_18\
        );

    \I__4255\ : InMux
    port map (
            O => \N__29066\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_1\
        );

    \I__4254\ : InMux
    port map (
            O => \N__29063\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_2\
        );

    \I__4253\ : InMux
    port map (
            O => \N__29060\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_3\
        );

    \I__4252\ : InMux
    port map (
            O => \N__29057\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_4\
        );

    \I__4251\ : InMux
    port map (
            O => \N__29054\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_5\
        );

    \I__4250\ : InMux
    port map (
            O => \N__29051\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_6\
        );

    \I__4249\ : InMux
    port map (
            O => \N__29048\,
            I => \bfn_10_3_0_\
        );

    \I__4248\ : InMux
    port map (
            O => \N__29045\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_8\
        );

    \I__4247\ : InMux
    port map (
            O => \N__29042\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_9\
        );

    \I__4246\ : InMux
    port map (
            O => \N__29039\,
            I => \N__29036\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__29036\,
            I => \N__29033\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__29033\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30\
        );

    \I__4243\ : InMux
    port map (
            O => \N__29030\,
            I => \N__29027\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__29027\,
            I => \N__29023\
        );

    \I__4241\ : CascadeMux
    port map (
            O => \N__29026\,
            I => \N__29020\
        );

    \I__4240\ : Span12Mux_s10_h
    port map (
            O => \N__29023\,
            I => \N__29016\
        );

    \I__4239\ : InMux
    port map (
            O => \N__29020\,
            I => \N__29011\
        );

    \I__4238\ : InMux
    port map (
            O => \N__29019\,
            I => \N__29011\
        );

    \I__4237\ : Span12Mux_v
    port map (
            O => \N__29016\,
            I => \N__29008\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__29011\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__4235\ : Odrv12
    port map (
            O => \N__29008\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__4234\ : IoInMux
    port map (
            O => \N__29003\,
            I => \N__29000\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__29000\,
            I => \N__28997\
        );

    \I__4232\ : Span4Mux_s3_v
    port map (
            O => \N__28997\,
            I => \N__28994\
        );

    \I__4231\ : Span4Mux_v
    port map (
            O => \N__28994\,
            I => \N__28991\
        );

    \I__4230\ : Odrv4
    port map (
            O => \N__28991\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__4229\ : InMux
    port map (
            O => \N__28988\,
            I => \N__28983\
        );

    \I__4228\ : InMux
    port map (
            O => \N__28987\,
            I => \N__28978\
        );

    \I__4227\ : InMux
    port map (
            O => \N__28986\,
            I => \N__28978\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__28983\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_30\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__28978\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_30\
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__28973\,
            I => \N__28969\
        );

    \I__4223\ : InMux
    port map (
            O => \N__28972\,
            I => \N__28962\
        );

    \I__4222\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28962\
        );

    \I__4221\ : InMux
    port map (
            O => \N__28968\,
            I => \N__28957\
        );

    \I__4220\ : InMux
    port map (
            O => \N__28967\,
            I => \N__28957\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__28962\,
            I => \N__28954\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__28957\,
            I => \N__28949\
        );

    \I__4217\ : Span12Mux_s8_v
    port map (
            O => \N__28954\,
            I => \N__28949\
        );

    \I__4216\ : Span12Mux_v
    port map (
            O => \N__28949\,
            I => \N__28946\
        );

    \I__4215\ : Odrv12
    port map (
            O => \N__28946\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28\
        );

    \I__4214\ : InMux
    port map (
            O => \N__28943\,
            I => \N__28938\
        );

    \I__4213\ : InMux
    port map (
            O => \N__28942\,
            I => \N__28933\
        );

    \I__4212\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28933\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__28938\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_31\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__28933\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_31\
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__28928\,
            I => \N__28925\
        );

    \I__4208\ : InMux
    port map (
            O => \N__28925\,
            I => \N__28922\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__28922\,
            I => \N__28919\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__28919\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt30\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__28916\,
            I => \N__28913\
        );

    \I__4204\ : InMux
    port map (
            O => \N__28913\,
            I => \N__28909\
        );

    \I__4203\ : InMux
    port map (
            O => \N__28912\,
            I => \N__28905\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__28909\,
            I => \N__28902\
        );

    \I__4201\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28899\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__28905\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_25\
        );

    \I__4199\ : Odrv4
    port map (
            O => \N__28902\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_25\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__28899\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_25\
        );

    \I__4197\ : InMux
    port map (
            O => \N__28892\,
            I => \N__28888\
        );

    \I__4196\ : InMux
    port map (
            O => \N__28891\,
            I => \N__28885\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__28888\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__28885\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__28880\,
            I => \N__28875\
        );

    \I__4192\ : InMux
    port map (
            O => \N__28879\,
            I => \N__28872\
        );

    \I__4191\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28867\
        );

    \I__4190\ : InMux
    port map (
            O => \N__28875\,
            I => \N__28867\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__28872\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_24\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__28867\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_24\
        );

    \I__4187\ : InMux
    port map (
            O => \N__28862\,
            I => \N__28856\
        );

    \I__4186\ : InMux
    port map (
            O => \N__28861\,
            I => \N__28856\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__28856\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_24\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__28853\,
            I => \N__28850\
        );

    \I__4183\ : InMux
    port map (
            O => \N__28850\,
            I => \N__28847\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__28847\,
            I => \N__28844\
        );

    \I__4181\ : Span4Mux_h
    port map (
            O => \N__28844\,
            I => \N__28841\
        );

    \I__4180\ : Odrv4
    port map (
            O => \N__28841\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt24\
        );

    \I__4179\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28818\
        );

    \I__4178\ : InMux
    port map (
            O => \N__28837\,
            I => \N__28818\
        );

    \I__4177\ : InMux
    port map (
            O => \N__28836\,
            I => \N__28818\
        );

    \I__4176\ : InMux
    port map (
            O => \N__28835\,
            I => \N__28818\
        );

    \I__4175\ : InMux
    port map (
            O => \N__28834\,
            I => \N__28797\
        );

    \I__4174\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28797\
        );

    \I__4173\ : InMux
    port map (
            O => \N__28832\,
            I => \N__28797\
        );

    \I__4172\ : InMux
    port map (
            O => \N__28831\,
            I => \N__28797\
        );

    \I__4171\ : InMux
    port map (
            O => \N__28830\,
            I => \N__28788\
        );

    \I__4170\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28788\
        );

    \I__4169\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28788\
        );

    \I__4168\ : InMux
    port map (
            O => \N__28827\,
            I => \N__28788\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__28818\,
            I => \N__28777\
        );

    \I__4166\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28768\
        );

    \I__4165\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28768\
        );

    \I__4164\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28768\
        );

    \I__4163\ : InMux
    port map (
            O => \N__28814\,
            I => \N__28768\
        );

    \I__4162\ : InMux
    port map (
            O => \N__28813\,
            I => \N__28759\
        );

    \I__4161\ : InMux
    port map (
            O => \N__28812\,
            I => \N__28759\
        );

    \I__4160\ : InMux
    port map (
            O => \N__28811\,
            I => \N__28759\
        );

    \I__4159\ : InMux
    port map (
            O => \N__28810\,
            I => \N__28759\
        );

    \I__4158\ : InMux
    port map (
            O => \N__28809\,
            I => \N__28750\
        );

    \I__4157\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28750\
        );

    \I__4156\ : InMux
    port map (
            O => \N__28807\,
            I => \N__28750\
        );

    \I__4155\ : InMux
    port map (
            O => \N__28806\,
            I => \N__28750\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__28797\,
            I => \N__28745\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__28788\,
            I => \N__28745\
        );

    \I__4152\ : InMux
    port map (
            O => \N__28787\,
            I => \N__28736\
        );

    \I__4151\ : InMux
    port map (
            O => \N__28786\,
            I => \N__28736\
        );

    \I__4150\ : InMux
    port map (
            O => \N__28785\,
            I => \N__28736\
        );

    \I__4149\ : InMux
    port map (
            O => \N__28784\,
            I => \N__28736\
        );

    \I__4148\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28727\
        );

    \I__4147\ : InMux
    port map (
            O => \N__28782\,
            I => \N__28727\
        );

    \I__4146\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28727\
        );

    \I__4145\ : InMux
    port map (
            O => \N__28780\,
            I => \N__28727\
        );

    \I__4144\ : Span4Mux_h
    port map (
            O => \N__28777\,
            I => \N__28722\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__28768\,
            I => \N__28722\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__28759\,
            I => \N__28715\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__28750\,
            I => \N__28715\
        );

    \I__4140\ : Span4Mux_h
    port map (
            O => \N__28745\,
            I => \N__28715\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__28736\,
            I => \phase_controller_inst1.stoper_tr.start_latched_i_0\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__28727\,
            I => \phase_controller_inst1.stoper_tr.start_latched_i_0\
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__28722\,
            I => \phase_controller_inst1.stoper_tr.start_latched_i_0\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__28715\,
            I => \phase_controller_inst1.stoper_tr.start_latched_i_0\
        );

    \I__4135\ : InMux
    port map (
            O => \N__28706\,
            I => \N__28703\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__28703\,
            I => \N__28700\
        );

    \I__4133\ : Span4Mux_h
    port map (
            O => \N__28700\,
            I => \N__28696\
        );

    \I__4132\ : CascadeMux
    port map (
            O => \N__28699\,
            I => \N__28692\
        );

    \I__4131\ : Sp12to4
    port map (
            O => \N__28696\,
            I => \N__28688\
        );

    \I__4130\ : InMux
    port map (
            O => \N__28695\,
            I => \N__28683\
        );

    \I__4129\ : InMux
    port map (
            O => \N__28692\,
            I => \N__28683\
        );

    \I__4128\ : InMux
    port map (
            O => \N__28691\,
            I => \N__28680\
        );

    \I__4127\ : Span12Mux_v
    port map (
            O => \N__28688\,
            I => \N__28677\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__28683\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__28680\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4124\ : Odrv12
    port map (
            O => \N__28677\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4123\ : IoInMux
    port map (
            O => \N__28670\,
            I => \N__28667\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__28667\,
            I => \N__28664\
        );

    \I__4121\ : Odrv4
    port map (
            O => \N__28664\,
            I => s3_phy_c
        );

    \I__4120\ : InMux
    port map (
            O => \N__28661\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_0\
        );

    \I__4119\ : InMux
    port map (
            O => \N__28658\,
            I => \N__28655\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__28655\,
            I => \N__28652\
        );

    \I__4117\ : Span4Mux_h
    port map (
            O => \N__28652\,
            I => \N__28648\
        );

    \I__4116\ : InMux
    port map (
            O => \N__28651\,
            I => \N__28645\
        );

    \I__4115\ : Odrv4
    port map (
            O => \N__28648\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__28645\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16\
        );

    \I__4113\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28635\
        );

    \I__4112\ : InMux
    port map (
            O => \N__28639\,
            I => \N__28632\
        );

    \I__4111\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28629\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__28635\,
            I => \N__28626\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__28632\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_17\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__28629\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_17\
        );

    \I__4107\ : Odrv4
    port map (
            O => \N__28626\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_17\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__28619\,
            I => \N__28615\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__28618\,
            I => \N__28611\
        );

    \I__4104\ : InMux
    port map (
            O => \N__28615\,
            I => \N__28608\
        );

    \I__4103\ : InMux
    port map (
            O => \N__28614\,
            I => \N__28605\
        );

    \I__4102\ : InMux
    port map (
            O => \N__28611\,
            I => \N__28602\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__28608\,
            I => \N__28599\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__28605\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_16\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__28602\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_16\
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__28599\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_16\
        );

    \I__4097\ : InMux
    port map (
            O => \N__28592\,
            I => \N__28589\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__28589\,
            I => \N__28586\
        );

    \I__4095\ : Span4Mux_h
    port map (
            O => \N__28586\,
            I => \N__28582\
        );

    \I__4094\ : InMux
    port map (
            O => \N__28585\,
            I => \N__28579\
        );

    \I__4093\ : Odrv4
    port map (
            O => \N__28582\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__28579\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17\
        );

    \I__4091\ : InMux
    port map (
            O => \N__28574\,
            I => \N__28571\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__28571\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt16\
        );

    \I__4089\ : InMux
    port map (
            O => \N__28568\,
            I => \N__28562\
        );

    \I__4088\ : InMux
    port map (
            O => \N__28567\,
            I => \N__28562\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__28562\,
            I => \N__28558\
        );

    \I__4086\ : InMux
    port map (
            O => \N__28561\,
            I => \N__28555\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__28558\,
            I => \N__28552\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__28555\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_28\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__28552\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_28\
        );

    \I__4082\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28540\
        );

    \I__4081\ : InMux
    port map (
            O => \N__28546\,
            I => \N__28540\
        );

    \I__4080\ : InMux
    port map (
            O => \N__28545\,
            I => \N__28537\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__28540\,
            I => \N__28534\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__28537\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_29\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__28534\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_29\
        );

    \I__4076\ : InMux
    port map (
            O => \N__28529\,
            I => \N__28526\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__28526\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt28\
        );

    \I__4074\ : InMux
    port map (
            O => \N__28523\,
            I => \N__28520\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__28520\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22\
        );

    \I__4072\ : InMux
    port map (
            O => \N__28517\,
            I => \N__28514\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__28514\,
            I => \N__28511\
        );

    \I__4070\ : Span4Mux_v
    port map (
            O => \N__28511\,
            I => \N__28507\
        );

    \I__4069\ : InMux
    port map (
            O => \N__28510\,
            I => \N__28504\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__28507\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_24
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__28504\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_24
        );

    \I__4066\ : InMux
    port map (
            O => \N__28499\,
            I => \N__28495\
        );

    \I__4065\ : InMux
    port map (
            O => \N__28498\,
            I => \N__28492\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__28495\,
            I => \N__28489\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__28492\,
            I => \N__28486\
        );

    \I__4062\ : Span4Mux_v
    port map (
            O => \N__28489\,
            I => \N__28481\
        );

    \I__4061\ : Span4Mux_v
    port map (
            O => \N__28486\,
            I => \N__28481\
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__28481\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_25
        );

    \I__4059\ : InMux
    port map (
            O => \N__28478\,
            I => \N__28475\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__28475\,
            I => \N__28472\
        );

    \I__4057\ : Odrv4
    port map (
            O => \N__28472\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt26\
        );

    \I__4056\ : InMux
    port map (
            O => \N__28469\,
            I => \N__28466\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__28466\,
            I => \N__28462\
        );

    \I__4054\ : InMux
    port map (
            O => \N__28465\,
            I => \N__28459\
        );

    \I__4053\ : Span4Mux_h
    port map (
            O => \N__28462\,
            I => \N__28456\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__28459\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_26
        );

    \I__4051\ : Odrv4
    port map (
            O => \N__28456\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_26
        );

    \I__4050\ : InMux
    port map (
            O => \N__28451\,
            I => \N__28446\
        );

    \I__4049\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28441\
        );

    \I__4048\ : InMux
    port map (
            O => \N__28449\,
            I => \N__28441\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__28446\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_27\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__28441\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_27\
        );

    \I__4045\ : InMux
    port map (
            O => \N__28436\,
            I => \N__28430\
        );

    \I__4044\ : InMux
    port map (
            O => \N__28435\,
            I => \N__28430\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__28430\,
            I => \N__28427\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__28427\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__28424\,
            I => \N__28420\
        );

    \I__4040\ : CascadeMux
    port map (
            O => \N__28423\,
            I => \N__28417\
        );

    \I__4039\ : InMux
    port map (
            O => \N__28420\,
            I => \N__28412\
        );

    \I__4038\ : InMux
    port map (
            O => \N__28417\,
            I => \N__28412\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__28412\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26\
        );

    \I__4036\ : InMux
    port map (
            O => \N__28409\,
            I => \N__28404\
        );

    \I__4035\ : InMux
    port map (
            O => \N__28408\,
            I => \N__28399\
        );

    \I__4034\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28399\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__28404\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_26\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__28399\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_26\
        );

    \I__4031\ : CascadeMux
    port map (
            O => \N__28394\,
            I => \N__28391\
        );

    \I__4030\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28388\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__28388\,
            I => \N__28385\
        );

    \I__4028\ : Odrv4
    port map (
            O => \N__28385\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26\
        );

    \I__4027\ : InMux
    port map (
            O => \N__28382\,
            I => \N__28379\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__28379\,
            I => \N__28376\
        );

    \I__4025\ : Odrv4
    port map (
            O => \N__28376\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24\
        );

    \I__4024\ : InMux
    port map (
            O => \N__28373\,
            I => \bfn_9_21_0_\
        );

    \I__4023\ : InMux
    port map (
            O => \N__28370\,
            I => \N__28364\
        );

    \I__4022\ : InMux
    port map (
            O => \N__28369\,
            I => \N__28364\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__28364\,
            I => \N__28360\
        );

    \I__4020\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28357\
        );

    \I__4019\ : Odrv12
    port map (
            O => \N__28360\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__28357\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__28352\,
            I => \N__28348\
        );

    \I__4016\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28345\
        );

    \I__4015\ : InMux
    port map (
            O => \N__28348\,
            I => \N__28342\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__28345\,
            I => \phase_controller_inst1.stoper_tr.counter\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__28342\,
            I => \phase_controller_inst1.stoper_tr.counter\
        );

    \I__4012\ : CascadeMux
    port map (
            O => \N__28337\,
            I => \N__28334\
        );

    \I__4011\ : InMux
    port map (
            O => \N__28334\,
            I => \N__28331\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__28331\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28\
        );

    \I__4009\ : InMux
    port map (
            O => \N__28328\,
            I => \N__28325\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__28325\,
            I => \N__28322\
        );

    \I__4007\ : Span4Mux_v
    port map (
            O => \N__28322\,
            I => \N__28319\
        );

    \I__4006\ : Odrv4
    port map (
            O => \N__28319\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_11\
        );

    \I__4005\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28312\
        );

    \I__4004\ : InMux
    port map (
            O => \N__28315\,
            I => \N__28309\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__28312\,
            I => \N__28306\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__28309\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_11\
        );

    \I__4001\ : Odrv4
    port map (
            O => \N__28306\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_11\
        );

    \I__4000\ : CascadeMux
    port map (
            O => \N__28301\,
            I => \N__28298\
        );

    \I__3999\ : InMux
    port map (
            O => \N__28298\,
            I => \N__28295\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__28295\,
            I => \phase_controller_inst1.stoper_tr.counter_i_11\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__28292\,
            I => \N__28289\
        );

    \I__3996\ : InMux
    port map (
            O => \N__28289\,
            I => \N__28286\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__28286\,
            I => \N__28283\
        );

    \I__3994\ : Span4Mux_v
    port map (
            O => \N__28283\,
            I => \N__28280\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__28280\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_12\
        );

    \I__3992\ : InMux
    port map (
            O => \N__28277\,
            I => \N__28273\
        );

    \I__3991\ : InMux
    port map (
            O => \N__28276\,
            I => \N__28270\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__28273\,
            I => \N__28267\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__28270\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_12\
        );

    \I__3988\ : Odrv4
    port map (
            O => \N__28267\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_12\
        );

    \I__3987\ : InMux
    port map (
            O => \N__28262\,
            I => \N__28259\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__28259\,
            I => \phase_controller_inst1.stoper_tr.counter_i_12\
        );

    \I__3985\ : InMux
    port map (
            O => \N__28256\,
            I => \N__28252\
        );

    \I__3984\ : InMux
    port map (
            O => \N__28255\,
            I => \N__28249\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__28252\,
            I => \N__28246\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__28249\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_13\
        );

    \I__3981\ : Odrv4
    port map (
            O => \N__28246\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_13\
        );

    \I__3980\ : InMux
    port map (
            O => \N__28241\,
            I => \N__28238\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__28238\,
            I => \N__28235\
        );

    \I__3978\ : Span4Mux_v
    port map (
            O => \N__28235\,
            I => \N__28232\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__28232\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_13\
        );

    \I__3976\ : CascadeMux
    port map (
            O => \N__28229\,
            I => \N__28226\
        );

    \I__3975\ : InMux
    port map (
            O => \N__28226\,
            I => \N__28223\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__28223\,
            I => \phase_controller_inst1.stoper_tr.counter_i_13\
        );

    \I__3973\ : InMux
    port map (
            O => \N__28220\,
            I => \N__28216\
        );

    \I__3972\ : InMux
    port map (
            O => \N__28219\,
            I => \N__28213\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__28216\,
            I => \N__28210\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__28213\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_14\
        );

    \I__3969\ : Odrv4
    port map (
            O => \N__28210\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_14\
        );

    \I__3968\ : InMux
    port map (
            O => \N__28205\,
            I => \N__28202\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__28202\,
            I => \N__28199\
        );

    \I__3966\ : Span4Mux_h
    port map (
            O => \N__28199\,
            I => \N__28196\
        );

    \I__3965\ : Odrv4
    port map (
            O => \N__28196\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_14\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__28193\,
            I => \N__28190\
        );

    \I__3963\ : InMux
    port map (
            O => \N__28190\,
            I => \N__28187\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__28187\,
            I => \phase_controller_inst1.stoper_tr.counter_i_14\
        );

    \I__3961\ : InMux
    port map (
            O => \N__28184\,
            I => \N__28180\
        );

    \I__3960\ : InMux
    port map (
            O => \N__28183\,
            I => \N__28177\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__28180\,
            I => \N__28174\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__28177\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_15\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__28174\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_15\
        );

    \I__3956\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28166\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__28166\,
            I => \N__28163\
        );

    \I__3954\ : Span4Mux_h
    port map (
            O => \N__28163\,
            I => \N__28160\
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__28160\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_15\
        );

    \I__3952\ : CascadeMux
    port map (
            O => \N__28157\,
            I => \N__28154\
        );

    \I__3951\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28151\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__28151\,
            I => \phase_controller_inst1.stoper_tr.counter_i_15\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__28148\,
            I => \N__28145\
        );

    \I__3948\ : InMux
    port map (
            O => \N__28145\,
            I => \N__28142\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__28142\,
            I => \N__28139\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__28139\,
            I => \N__28136\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__28136\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16\
        );

    \I__3944\ : InMux
    port map (
            O => \N__28133\,
            I => \N__28130\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__28130\,
            I => \N__28127\
        );

    \I__3942\ : Odrv12
    port map (
            O => \N__28127\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__28124\,
            I => \N__28121\
        );

    \I__3940\ : InMux
    port map (
            O => \N__28121\,
            I => \N__28118\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__28118\,
            I => \N__28115\
        );

    \I__3938\ : Odrv4
    port map (
            O => \N__28115\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt18\
        );

    \I__3937\ : CascadeMux
    port map (
            O => \N__28112\,
            I => \N__28109\
        );

    \I__3936\ : InMux
    port map (
            O => \N__28109\,
            I => \N__28106\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__28106\,
            I => \phase_controller_inst1.stoper_tr.counter_i_3\
        );

    \I__3934\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28100\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__28100\,
            I => \N__28097\
        );

    \I__3932\ : Odrv12
    port map (
            O => \N__28097\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_4\
        );

    \I__3931\ : InMux
    port map (
            O => \N__28094\,
            I => \N__28090\
        );

    \I__3930\ : InMux
    port map (
            O => \N__28093\,
            I => \N__28087\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__28090\,
            I => \N__28084\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__28087\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_4\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__28084\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_4\
        );

    \I__3926\ : CascadeMux
    port map (
            O => \N__28079\,
            I => \N__28076\
        );

    \I__3925\ : InMux
    port map (
            O => \N__28076\,
            I => \N__28073\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__28073\,
            I => \N__28070\
        );

    \I__3923\ : Odrv4
    port map (
            O => \N__28070\,
            I => \phase_controller_inst1.stoper_tr.counter_i_4\
        );

    \I__3922\ : InMux
    port map (
            O => \N__28067\,
            I => \N__28063\
        );

    \I__3921\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28060\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__28063\,
            I => \N__28057\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__28060\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_5\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__28057\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_5\
        );

    \I__3917\ : InMux
    port map (
            O => \N__28052\,
            I => \N__28049\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__28049\,
            I => \N__28046\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__28046\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_5\
        );

    \I__3914\ : CascadeMux
    port map (
            O => \N__28043\,
            I => \N__28040\
        );

    \I__3913\ : InMux
    port map (
            O => \N__28040\,
            I => \N__28037\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__28037\,
            I => \phase_controller_inst1.stoper_tr.counter_i_5\
        );

    \I__3911\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28030\
        );

    \I__3910\ : InMux
    port map (
            O => \N__28033\,
            I => \N__28027\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__28030\,
            I => \N__28024\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__28027\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_6\
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__28024\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_6\
        );

    \I__3906\ : InMux
    port map (
            O => \N__28019\,
            I => \N__28016\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__28016\,
            I => \N__28013\
        );

    \I__3904\ : Odrv12
    port map (
            O => \N__28013\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_6\
        );

    \I__3903\ : CascadeMux
    port map (
            O => \N__28010\,
            I => \N__28007\
        );

    \I__3902\ : InMux
    port map (
            O => \N__28007\,
            I => \N__28004\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__28004\,
            I => \phase_controller_inst1.stoper_tr.counter_i_6\
        );

    \I__3900\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27998\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__27998\,
            I => \N__27994\
        );

    \I__3898\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27991\
        );

    \I__3897\ : Span4Mux_v
    port map (
            O => \N__27994\,
            I => \N__27988\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__27991\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_7\
        );

    \I__3895\ : Odrv4
    port map (
            O => \N__27988\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_7\
        );

    \I__3894\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27980\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__27980\,
            I => \N__27977\
        );

    \I__3892\ : Odrv4
    port map (
            O => \N__27977\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_7\
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__27974\,
            I => \N__27971\
        );

    \I__3890\ : InMux
    port map (
            O => \N__27971\,
            I => \N__27968\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__27968\,
            I => \phase_controller_inst1.stoper_tr.counter_i_7\
        );

    \I__3888\ : CascadeMux
    port map (
            O => \N__27965\,
            I => \N__27962\
        );

    \I__3887\ : InMux
    port map (
            O => \N__27962\,
            I => \N__27959\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__27959\,
            I => \N__27956\
        );

    \I__3885\ : Span4Mux_v
    port map (
            O => \N__27956\,
            I => \N__27953\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__27953\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_8\
        );

    \I__3883\ : InMux
    port map (
            O => \N__27950\,
            I => \N__27947\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__27947\,
            I => \N__27943\
        );

    \I__3881\ : InMux
    port map (
            O => \N__27946\,
            I => \N__27940\
        );

    \I__3880\ : Span4Mux_h
    port map (
            O => \N__27943\,
            I => \N__27937\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__27940\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_8\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__27937\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_8\
        );

    \I__3877\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27929\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__27929\,
            I => \phase_controller_inst1.stoper_tr.counter_i_8\
        );

    \I__3875\ : InMux
    port map (
            O => \N__27926\,
            I => \N__27923\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__27923\,
            I => \N__27920\
        );

    \I__3873\ : Span4Mux_v
    port map (
            O => \N__27920\,
            I => \N__27917\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__27917\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_9\
        );

    \I__3871\ : InMux
    port map (
            O => \N__27914\,
            I => \N__27910\
        );

    \I__3870\ : InMux
    port map (
            O => \N__27913\,
            I => \N__27907\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__27910\,
            I => \N__27904\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__27907\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_9\
        );

    \I__3867\ : Odrv4
    port map (
            O => \N__27904\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_9\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__27899\,
            I => \N__27896\
        );

    \I__3865\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27893\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__27893\,
            I => \phase_controller_inst1.stoper_tr.counter_i_9\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__27890\,
            I => \N__27887\
        );

    \I__3862\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27884\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__27884\,
            I => \N__27881\
        );

    \I__3860\ : Span4Mux_v
    port map (
            O => \N__27881\,
            I => \N__27878\
        );

    \I__3859\ : Odrv4
    port map (
            O => \N__27878\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_10\
        );

    \I__3858\ : InMux
    port map (
            O => \N__27875\,
            I => \N__27871\
        );

    \I__3857\ : InMux
    port map (
            O => \N__27874\,
            I => \N__27868\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__27871\,
            I => \N__27865\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__27868\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_10\
        );

    \I__3854\ : Odrv4
    port map (
            O => \N__27865\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_10\
        );

    \I__3853\ : InMux
    port map (
            O => \N__27860\,
            I => \N__27857\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__27857\,
            I => \phase_controller_inst1.stoper_tr.counter_i_10\
        );

    \I__3851\ : InMux
    port map (
            O => \N__27854\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27\
        );

    \I__3850\ : InMux
    port map (
            O => \N__27851\,
            I => \N__27848\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__27848\,
            I => \N__27844\
        );

    \I__3848\ : InMux
    port map (
            O => \N__27847\,
            I => \N__27841\
        );

    \I__3847\ : Span4Mux_h
    port map (
            O => \N__27844\,
            I => \N__27838\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__27841\,
            I => \N__27835\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__27838\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__27835\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0\
        );

    \I__3843\ : InMux
    port map (
            O => \N__27830\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28\
        );

    \I__3842\ : InMux
    port map (
            O => \N__27827\,
            I => \N__27823\
        );

    \I__3841\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27820\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__27823\,
            I => \N__27817\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__27820\,
            I => \N__27812\
        );

    \I__3838\ : Span4Mux_h
    port map (
            O => \N__27817\,
            I => \N__27812\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__27812\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0\
        );

    \I__3836\ : InMux
    port map (
            O => \N__27809\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29\
        );

    \I__3835\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27803\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__27803\,
            I => \N__27800\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__27800\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO\
        );

    \I__3832\ : InMux
    port map (
            O => \N__27797\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30\
        );

    \I__3831\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27790\
        );

    \I__3830\ : InMux
    port map (
            O => \N__27793\,
            I => \N__27787\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__27790\,
            I => \N__27784\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__27787\,
            I => \N__27781\
        );

    \I__3827\ : Span4Mux_v
    port map (
            O => \N__27784\,
            I => \N__27778\
        );

    \I__3826\ : Span4Mux_h
    port map (
            O => \N__27781\,
            I => \N__27775\
        );

    \I__3825\ : Span4Mux_v
    port map (
            O => \N__27778\,
            I => \N__27772\
        );

    \I__3824\ : Odrv4
    port map (
            O => \N__27775\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_28
        );

    \I__3823\ : Odrv4
    port map (
            O => \N__27772\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_28
        );

    \I__3822\ : InMux
    port map (
            O => \N__27767\,
            I => \N__27764\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__27764\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29\
        );

    \I__3820\ : InMux
    port map (
            O => \N__27761\,
            I => \N__27758\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__27758\,
            I => \N__27754\
        );

    \I__3818\ : InMux
    port map (
            O => \N__27757\,
            I => \N__27751\
        );

    \I__3817\ : Span4Mux_h
    port map (
            O => \N__27754\,
            I => \N__27748\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__27751\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_0\
        );

    \I__3815\ : Odrv4
    port map (
            O => \N__27748\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_0\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__27743\,
            I => \N__27740\
        );

    \I__3813\ : InMux
    port map (
            O => \N__27740\,
            I => \N__27737\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__27737\,
            I => \phase_controller_inst1.stoper_tr.counter_i_0\
        );

    \I__3811\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27731\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__27731\,
            I => \N__27728\
        );

    \I__3809\ : Span4Mux_v
    port map (
            O => \N__27728\,
            I => \N__27725\
        );

    \I__3808\ : Odrv4
    port map (
            O => \N__27725\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ1Z_1\
        );

    \I__3807\ : InMux
    port map (
            O => \N__27722\,
            I => \N__27718\
        );

    \I__3806\ : InMux
    port map (
            O => \N__27721\,
            I => \N__27715\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__27718\,
            I => \N__27712\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__27715\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_1\
        );

    \I__3803\ : Odrv4
    port map (
            O => \N__27712\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_1\
        );

    \I__3802\ : CascadeMux
    port map (
            O => \N__27707\,
            I => \N__27704\
        );

    \I__3801\ : InMux
    port map (
            O => \N__27704\,
            I => \N__27701\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__27701\,
            I => \N__27698\
        );

    \I__3799\ : Odrv4
    port map (
            O => \N__27698\,
            I => \phase_controller_inst1.stoper_tr.counter_i_1\
        );

    \I__3798\ : InMux
    port map (
            O => \N__27695\,
            I => \N__27692\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__27692\,
            I => \N__27689\
        );

    \I__3796\ : Span4Mux_h
    port map (
            O => \N__27689\,
            I => \N__27686\
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__27686\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_2\
        );

    \I__3794\ : InMux
    port map (
            O => \N__27683\,
            I => \N__27679\
        );

    \I__3793\ : InMux
    port map (
            O => \N__27682\,
            I => \N__27676\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__27679\,
            I => \N__27673\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__27676\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_2\
        );

    \I__3790\ : Odrv4
    port map (
            O => \N__27673\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_2\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__27668\,
            I => \N__27665\
        );

    \I__3788\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27662\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__27662\,
            I => \phase_controller_inst1.stoper_tr.counter_i_2\
        );

    \I__3786\ : InMux
    port map (
            O => \N__27659\,
            I => \N__27656\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__27656\,
            I => \N__27653\
        );

    \I__3784\ : Span4Mux_h
    port map (
            O => \N__27653\,
            I => \N__27650\
        );

    \I__3783\ : Odrv4
    port map (
            O => \N__27650\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_3\
        );

    \I__3782\ : InMux
    port map (
            O => \N__27647\,
            I => \N__27643\
        );

    \I__3781\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27640\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__27643\,
            I => \N__27637\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__27640\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_3\
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__27637\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_3\
        );

    \I__3777\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27629\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__27629\,
            I => \N__27625\
        );

    \I__3775\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27622\
        );

    \I__3774\ : Span4Mux_v
    port map (
            O => \N__27625\,
            I => \N__27619\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__27622\,
            I => \N__27616\
        );

    \I__3772\ : Odrv4
    port map (
            O => \N__27619\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__27616\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0\
        );

    \I__3770\ : InMux
    port map (
            O => \N__27611\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19\
        );

    \I__3769\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27605\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__27605\,
            I => \N__27602\
        );

    \I__3767\ : Odrv12
    port map (
            O => \N__27602\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21\
        );

    \I__3766\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27596\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__27596\,
            I => \N__27592\
        );

    \I__3764\ : InMux
    port map (
            O => \N__27595\,
            I => \N__27589\
        );

    \I__3763\ : Span4Mux_h
    port map (
            O => \N__27592\,
            I => \N__27586\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__27589\,
            I => \N__27583\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__27586\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__27583\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0\
        );

    \I__3759\ : InMux
    port map (
            O => \N__27578\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20\
        );

    \I__3758\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27571\
        );

    \I__3757\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27568\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__27571\,
            I => \N__27565\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__27568\,
            I => \N__27560\
        );

    \I__3754\ : Span4Mux_h
    port map (
            O => \N__27565\,
            I => \N__27560\
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__27560\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0\
        );

    \I__3752\ : InMux
    port map (
            O => \N__27557\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21\
        );

    \I__3751\ : InMux
    port map (
            O => \N__27554\,
            I => \N__27551\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__27551\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23\
        );

    \I__3749\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27545\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__27545\,
            I => \N__27541\
        );

    \I__3747\ : InMux
    port map (
            O => \N__27544\,
            I => \N__27538\
        );

    \I__3746\ : Span4Mux_h
    port map (
            O => \N__27541\,
            I => \N__27533\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__27538\,
            I => \N__27533\
        );

    \I__3744\ : Odrv4
    port map (
            O => \N__27533\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0\
        );

    \I__3743\ : InMux
    port map (
            O => \N__27530\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22\
        );

    \I__3742\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27523\
        );

    \I__3741\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27520\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__27523\,
            I => \N__27517\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__27520\,
            I => \N__27512\
        );

    \I__3738\ : Span4Mux_h
    port map (
            O => \N__27517\,
            I => \N__27512\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__27512\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0\
        );

    \I__3736\ : InMux
    port map (
            O => \N__27509\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23\
        );

    \I__3735\ : InMux
    port map (
            O => \N__27506\,
            I => \N__27502\
        );

    \I__3734\ : InMux
    port map (
            O => \N__27505\,
            I => \N__27499\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__27502\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__27499\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0\
        );

    \I__3731\ : InMux
    port map (
            O => \N__27494\,
            I => \bfn_9_17_0_\
        );

    \I__3730\ : InMux
    port map (
            O => \N__27491\,
            I => \N__27487\
        );

    \I__3729\ : InMux
    port map (
            O => \N__27490\,
            I => \N__27484\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__27487\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__27484\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0\
        );

    \I__3726\ : InMux
    port map (
            O => \N__27479\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25\
        );

    \I__3725\ : InMux
    port map (
            O => \N__27476\,
            I => \N__27472\
        );

    \I__3724\ : InMux
    port map (
            O => \N__27475\,
            I => \N__27469\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__27472\,
            I => \N__27464\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__27469\,
            I => \N__27464\
        );

    \I__3721\ : Span4Mux_v
    port map (
            O => \N__27464\,
            I => \N__27461\
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__27461\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0\
        );

    \I__3719\ : InMux
    port map (
            O => \N__27458\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26\
        );

    \I__3718\ : InMux
    port map (
            O => \N__27455\,
            I => \N__27452\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__27452\,
            I => \N__27448\
        );

    \I__3716\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27445\
        );

    \I__3715\ : Span4Mux_v
    port map (
            O => \N__27448\,
            I => \N__27442\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__27445\,
            I => \N__27439\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__27442\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0\
        );

    \I__3712\ : Odrv4
    port map (
            O => \N__27439\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0\
        );

    \I__3711\ : InMux
    port map (
            O => \N__27434\,
            I => \N__27431\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__27431\,
            I => \N__27427\
        );

    \I__3709\ : InMux
    port map (
            O => \N__27430\,
            I => \N__27424\
        );

    \I__3708\ : Span4Mux_v
    port map (
            O => \N__27427\,
            I => \N__27421\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__27424\,
            I => \N__27418\
        );

    \I__3706\ : Odrv4
    port map (
            O => \N__27421\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9\
        );

    \I__3705\ : Odrv4
    port map (
            O => \N__27418\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9\
        );

    \I__3704\ : InMux
    port map (
            O => \N__27413\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11\
        );

    \I__3703\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27407\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__27407\,
            I => \N__27403\
        );

    \I__3701\ : InMux
    port map (
            O => \N__27406\,
            I => \N__27400\
        );

    \I__3700\ : Span4Mux_h
    port map (
            O => \N__27403\,
            I => \N__27397\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__27400\,
            I => \N__27394\
        );

    \I__3698\ : Odrv4
    port map (
            O => \N__27397\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9\
        );

    \I__3697\ : Odrv4
    port map (
            O => \N__27394\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9\
        );

    \I__3696\ : InMux
    port map (
            O => \N__27389\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12\
        );

    \I__3695\ : InMux
    port map (
            O => \N__27386\,
            I => \N__27383\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__27383\,
            I => \N__27380\
        );

    \I__3693\ : Span4Mux_v
    port map (
            O => \N__27380\,
            I => \N__27377\
        );

    \I__3692\ : Odrv4
    port map (
            O => \N__27377\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14\
        );

    \I__3691\ : InMux
    port map (
            O => \N__27374\,
            I => \N__27370\
        );

    \I__3690\ : InMux
    port map (
            O => \N__27373\,
            I => \N__27367\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__27370\,
            I => \N__27364\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__27367\,
            I => \N__27359\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__27364\,
            I => \N__27359\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__27359\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9\
        );

    \I__3685\ : InMux
    port map (
            O => \N__27356\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13\
        );

    \I__3684\ : CascadeMux
    port map (
            O => \N__27353\,
            I => \N__27350\
        );

    \I__3683\ : InMux
    port map (
            O => \N__27350\,
            I => \N__27347\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__27347\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15\
        );

    \I__3681\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27341\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__27341\,
            I => \N__27337\
        );

    \I__3679\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27334\
        );

    \I__3678\ : Span4Mux_h
    port map (
            O => \N__27337\,
            I => \N__27331\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__27334\,
            I => \N__27328\
        );

    \I__3676\ : Odrv4
    port map (
            O => \N__27331\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9\
        );

    \I__3675\ : Odrv4
    port map (
            O => \N__27328\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9\
        );

    \I__3674\ : InMux
    port map (
            O => \N__27323\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14\
        );

    \I__3673\ : InMux
    port map (
            O => \N__27320\,
            I => \N__27316\
        );

    \I__3672\ : InMux
    port map (
            O => \N__27319\,
            I => \N__27313\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__27316\,
            I => \N__27310\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__27313\,
            I => \N__27305\
        );

    \I__3669\ : Span4Mux_h
    port map (
            O => \N__27310\,
            I => \N__27305\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__27305\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9\
        );

    \I__3667\ : InMux
    port map (
            O => \N__27302\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15\
        );

    \I__3666\ : InMux
    port map (
            O => \N__27299\,
            I => \N__27295\
        );

    \I__3665\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27292\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__27295\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__27292\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0\
        );

    \I__3662\ : InMux
    port map (
            O => \N__27287\,
            I => \bfn_9_16_0_\
        );

    \I__3661\ : InMux
    port map (
            O => \N__27284\,
            I => \N__27280\
        );

    \I__3660\ : InMux
    port map (
            O => \N__27283\,
            I => \N__27277\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__27280\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__27277\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0\
        );

    \I__3657\ : InMux
    port map (
            O => \N__27272\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17\
        );

    \I__3656\ : InMux
    port map (
            O => \N__27269\,
            I => \N__27265\
        );

    \I__3655\ : InMux
    port map (
            O => \N__27268\,
            I => \N__27262\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__27265\,
            I => \N__27259\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__27262\,
            I => \N__27256\
        );

    \I__3652\ : Span4Mux_v
    port map (
            O => \N__27259\,
            I => \N__27253\
        );

    \I__3651\ : Odrv4
    port map (
            O => \N__27256\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0\
        );

    \I__3650\ : Odrv4
    port map (
            O => \N__27253\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0\
        );

    \I__3649\ : InMux
    port map (
            O => \N__27248\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18\
        );

    \I__3648\ : InMux
    port map (
            O => \N__27245\,
            I => \N__27242\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__27242\,
            I => \N__27238\
        );

    \I__3646\ : InMux
    port map (
            O => \N__27241\,
            I => \N__27235\
        );

    \I__3645\ : Span4Mux_v
    port map (
            O => \N__27238\,
            I => \N__27232\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__27235\,
            I => \N__27229\
        );

    \I__3643\ : Odrv4
    port map (
            O => \N__27232\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0\
        );

    \I__3642\ : Odrv4
    port map (
            O => \N__27229\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0\
        );

    \I__3641\ : InMux
    port map (
            O => \N__27224\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3\
        );

    \I__3640\ : InMux
    port map (
            O => \N__27221\,
            I => \N__27217\
        );

    \I__3639\ : InMux
    port map (
            O => \N__27220\,
            I => \N__27214\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__27217\,
            I => \N__27209\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__27214\,
            I => \N__27209\
        );

    \I__3636\ : Span4Mux_h
    port map (
            O => \N__27209\,
            I => \N__27206\
        );

    \I__3635\ : Odrv4
    port map (
            O => \N__27206\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0\
        );

    \I__3634\ : InMux
    port map (
            O => \N__27203\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4\
        );

    \I__3633\ : InMux
    port map (
            O => \N__27200\,
            I => \N__27196\
        );

    \I__3632\ : InMux
    port map (
            O => \N__27199\,
            I => \N__27193\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__27196\,
            I => \N__27190\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__27193\,
            I => \N__27185\
        );

    \I__3629\ : Span4Mux_h
    port map (
            O => \N__27190\,
            I => \N__27185\
        );

    \I__3628\ : Odrv4
    port map (
            O => \N__27185\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0\
        );

    \I__3627\ : InMux
    port map (
            O => \N__27182\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5\
        );

    \I__3626\ : InMux
    port map (
            O => \N__27179\,
            I => \N__27176\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__27176\,
            I => \N__27173\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__27173\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7\
        );

    \I__3623\ : InMux
    port map (
            O => \N__27170\,
            I => \N__27167\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__27167\,
            I => \N__27163\
        );

    \I__3621\ : InMux
    port map (
            O => \N__27166\,
            I => \N__27160\
        );

    \I__3620\ : Span4Mux_h
    port map (
            O => \N__27163\,
            I => \N__27157\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__27160\,
            I => \N__27154\
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__27157\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0\
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__27154\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0\
        );

    \I__3616\ : InMux
    port map (
            O => \N__27149\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6\
        );

    \I__3615\ : InMux
    port map (
            O => \N__27146\,
            I => \N__27142\
        );

    \I__3614\ : InMux
    port map (
            O => \N__27145\,
            I => \N__27139\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__27142\,
            I => \N__27136\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__27139\,
            I => \N__27131\
        );

    \I__3611\ : Span4Mux_h
    port map (
            O => \N__27136\,
            I => \N__27131\
        );

    \I__3610\ : Odrv4
    port map (
            O => \N__27131\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0\
        );

    \I__3609\ : InMux
    port map (
            O => \N__27128\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7\
        );

    \I__3608\ : InMux
    port map (
            O => \N__27125\,
            I => \N__27121\
        );

    \I__3607\ : InMux
    port map (
            O => \N__27124\,
            I => \N__27118\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__27121\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__27118\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0\
        );

    \I__3604\ : InMux
    port map (
            O => \N__27113\,
            I => \bfn_9_15_0_\
        );

    \I__3603\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27106\
        );

    \I__3602\ : InMux
    port map (
            O => \N__27109\,
            I => \N__27103\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__27106\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__27103\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0\
        );

    \I__3599\ : InMux
    port map (
            O => \N__27098\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9\
        );

    \I__3598\ : InMux
    port map (
            O => \N__27095\,
            I => \N__27091\
        );

    \I__3597\ : InMux
    port map (
            O => \N__27094\,
            I => \N__27088\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__27091\,
            I => \N__27083\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__27088\,
            I => \N__27083\
        );

    \I__3594\ : Span4Mux_v
    port map (
            O => \N__27083\,
            I => \N__27080\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__27080\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9\
        );

    \I__3592\ : InMux
    port map (
            O => \N__27077\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10\
        );

    \I__3591\ : InMux
    port map (
            O => \N__27074\,
            I => \N__27068\
        );

    \I__3590\ : InMux
    port map (
            O => \N__27073\,
            I => \N__27068\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__27068\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__3588\ : InMux
    port map (
            O => \N__27065\,
            I => \N__27059\
        );

    \I__3587\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27059\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__27059\,
            I => \N__27056\
        );

    \I__3585\ : Odrv4
    port map (
            O => \N__27056\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__3584\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27050\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__27050\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__27047\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3_cascade_\
        );

    \I__3581\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27040\
        );

    \I__3580\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27037\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__27040\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__27037\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__3577\ : CascadeMux
    port map (
            O => \N__27032\,
            I => \N__27029\
        );

    \I__3576\ : InMux
    port map (
            O => \N__27029\,
            I => \N__27026\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__27026\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1\
        );

    \I__3574\ : InMux
    port map (
            O => \N__27023\,
            I => \N__27019\
        );

    \I__3573\ : InMux
    port map (
            O => \N__27022\,
            I => \N__27016\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__27019\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__27016\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__3570\ : InMux
    port map (
            O => \N__27011\,
            I => \N__27008\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__27008\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2\
        );

    \I__3568\ : InMux
    port map (
            O => \N__27005\,
            I => \N__27002\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__27002\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3\
        );

    \I__3566\ : InMux
    port map (
            O => \N__26999\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2\
        );

    \I__3565\ : InMux
    port map (
            O => \N__26996\,
            I => \N__26993\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__26993\,
            I => \N__26989\
        );

    \I__3563\ : InMux
    port map (
            O => \N__26992\,
            I => \N__26986\
        );

    \I__3562\ : Span4Mux_s1_v
    port map (
            O => \N__26989\,
            I => \N__26981\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__26986\,
            I => \N__26981\
        );

    \I__3560\ : Span4Mux_v
    port map (
            O => \N__26981\,
            I => \N__26977\
        );

    \I__3559\ : InMux
    port map (
            O => \N__26980\,
            I => \N__26972\
        );

    \I__3558\ : Span4Mux_h
    port map (
            O => \N__26977\,
            I => \N__26966\
        );

    \I__3557\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26961\
        );

    \I__3556\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26961\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__26972\,
            I => \N__26958\
        );

    \I__3554\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26951\
        );

    \I__3553\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26951\
        );

    \I__3552\ : InMux
    port map (
            O => \N__26969\,
            I => \N__26951\
        );

    \I__3551\ : Sp12to4
    port map (
            O => \N__26966\,
            I => \N__26948\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__26961\,
            I => \N__26945\
        );

    \I__3549\ : Span4Mux_v
    port map (
            O => \N__26958\,
            I => \N__26940\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__26951\,
            I => \N__26940\
        );

    \I__3547\ : Span12Mux_s11_v
    port map (
            O => \N__26948\,
            I => \N__26937\
        );

    \I__3546\ : Span4Mux_v
    port map (
            O => \N__26945\,
            I => \N__26934\
        );

    \I__3545\ : Span4Mux_v
    port map (
            O => \N__26940\,
            I => \N__26931\
        );

    \I__3544\ : Span12Mux_v
    port map (
            O => \N__26937\,
            I => \N__26924\
        );

    \I__3543\ : Sp12to4
    port map (
            O => \N__26934\,
            I => \N__26924\
        );

    \I__3542\ : Sp12to4
    port map (
            O => \N__26931\,
            I => \N__26924\
        );

    \I__3541\ : Span12Mux_h
    port map (
            O => \N__26924\,
            I => \N__26921\
        );

    \I__3540\ : Odrv12
    port map (
            O => \N__26921\,
            I => start_stop_c
        );

    \I__3539\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26914\
        );

    \I__3538\ : CascadeMux
    port map (
            O => \N__26917\,
            I => \N__26911\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__26914\,
            I => \N__26907\
        );

    \I__3536\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26902\
        );

    \I__3535\ : InMux
    port map (
            O => \N__26910\,
            I => \N__26902\
        );

    \I__3534\ : Span4Mux_h
    port map (
            O => \N__26907\,
            I => \N__26899\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__26902\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__26899\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__26894\,
            I => \phase_controller_inst1.state_ns_0_0_1_cascade_\
        );

    \I__3530\ : InMux
    port map (
            O => \N__26891\,
            I => \N__26888\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__26888\,
            I => \N__26885\
        );

    \I__3528\ : Span4Mux_h
    port map (
            O => \N__26885\,
            I => \N__26880\
        );

    \I__3527\ : InMux
    port map (
            O => \N__26884\,
            I => \N__26875\
        );

    \I__3526\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26875\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__26880\,
            I => \phase_controller_inst1.start_flagZ0\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__26875\,
            I => \phase_controller_inst1.start_flagZ0\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__26870\,
            I => \phase_controller_inst1.stoper_tr.un4_start_0_cascade_\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__26867\,
            I => \N__26862\
        );

    \I__3521\ : InMux
    port map (
            O => \N__26866\,
            I => \N__26855\
        );

    \I__3520\ : InMux
    port map (
            O => \N__26865\,
            I => \N__26855\
        );

    \I__3519\ : InMux
    port map (
            O => \N__26862\,
            I => \N__26855\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__26855\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__3517\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26846\
        );

    \I__3516\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26846\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__26846\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__3514\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26840\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__26840\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__26837\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7_cascade_\
        );

    \I__3511\ : InMux
    port map (
            O => \N__26834\,
            I => \N__26830\
        );

    \I__3510\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26827\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__26830\,
            I => \N__26824\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__26827\,
            I => \N__26821\
        );

    \I__3507\ : Span4Mux_h
    port map (
            O => \N__26824\,
            I => \N__26817\
        );

    \I__3506\ : Span4Mux_h
    port map (
            O => \N__26821\,
            I => \N__26814\
        );

    \I__3505\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26811\
        );

    \I__3504\ : Span4Mux_v
    port map (
            O => \N__26817\,
            I => \N__26808\
        );

    \I__3503\ : Sp12to4
    port map (
            O => \N__26814\,
            I => \N__26803\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__26811\,
            I => \N__26803\
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__26808\,
            I => il_min_comp2_c
        );

    \I__3500\ : Odrv12
    port map (
            O => \N__26803\,
            I => il_min_comp2_c
        );

    \I__3499\ : InMux
    port map (
            O => \N__26798\,
            I => \N__26794\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__26797\,
            I => \N__26791\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__26794\,
            I => \N__26788\
        );

    \I__3496\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26783\
        );

    \I__3495\ : Sp12to4
    port map (
            O => \N__26788\,
            I => \N__26780\
        );

    \I__3494\ : InMux
    port map (
            O => \N__26787\,
            I => \N__26777\
        );

    \I__3493\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26774\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__26783\,
            I => \N__26771\
        );

    \I__3491\ : Span12Mux_v
    port map (
            O => \N__26780\,
            I => \N__26768\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__26777\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__26774\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3488\ : Odrv4
    port map (
            O => \N__26771\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3487\ : Odrv12
    port map (
            O => \N__26768\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3486\ : InMux
    port map (
            O => \N__26759\,
            I => \N__26753\
        );

    \I__3485\ : InMux
    port map (
            O => \N__26758\,
            I => \N__26753\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__26753\,
            I => \N__26749\
        );

    \I__3483\ : InMux
    port map (
            O => \N__26752\,
            I => \N__26746\
        );

    \I__3482\ : Span4Mux_v
    port map (
            O => \N__26749\,
            I => \N__26741\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__26746\,
            I => \N__26741\
        );

    \I__3480\ : Span4Mux_v
    port map (
            O => \N__26741\,
            I => \N__26738\
        );

    \I__3479\ : Span4Mux_h
    port map (
            O => \N__26738\,
            I => \N__26735\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__26735\,
            I => il_max_comp2_c
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__26732\,
            I => \N__26727\
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__26731\,
            I => \N__26724\
        );

    \I__3475\ : InMux
    port map (
            O => \N__26730\,
            I => \N__26716\
        );

    \I__3474\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26716\
        );

    \I__3473\ : InMux
    port map (
            O => \N__26724\,
            I => \N__26716\
        );

    \I__3472\ : InMux
    port map (
            O => \N__26723\,
            I => \N__26713\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__26716\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__26713\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__3469\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26699\
        );

    \I__3468\ : InMux
    port map (
            O => \N__26707\,
            I => \N__26699\
        );

    \I__3467\ : InMux
    port map (
            O => \N__26706\,
            I => \N__26691\
        );

    \I__3466\ : InMux
    port map (
            O => \N__26705\,
            I => \N__26691\
        );

    \I__3465\ : InMux
    port map (
            O => \N__26704\,
            I => \N__26691\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__26699\,
            I => \N__26688\
        );

    \I__3463\ : InMux
    port map (
            O => \N__26698\,
            I => \N__26685\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__26691\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__26688\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__26685\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__3459\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26673\
        );

    \I__3458\ : InMux
    port map (
            O => \N__26677\,
            I => \N__26668\
        );

    \I__3457\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26668\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__26673\,
            I => \N__26665\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__26668\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__3454\ : Odrv4
    port map (
            O => \N__26665\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__3453\ : InMux
    port map (
            O => \N__26660\,
            I => \N__26657\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__26657\,
            I => \phase_controller_inst2.stoper_hc.un4_start_0\
        );

    \I__3451\ : InMux
    port map (
            O => \N__26654\,
            I => \N__26644\
        );

    \I__3450\ : InMux
    port map (
            O => \N__26653\,
            I => \N__26644\
        );

    \I__3449\ : InMux
    port map (
            O => \N__26652\,
            I => \N__26644\
        );

    \I__3448\ : InMux
    port map (
            O => \N__26651\,
            I => \N__26641\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__26644\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__26641\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__3445\ : InMux
    port map (
            O => \N__26636\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_28\
        );

    \I__3444\ : InMux
    port map (
            O => \N__26633\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_29\
        );

    \I__3443\ : InMux
    port map (
            O => \N__26630\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_30\
        );

    \I__3442\ : CEMux
    port map (
            O => \N__26627\,
            I => \N__26615\
        );

    \I__3441\ : CEMux
    port map (
            O => \N__26626\,
            I => \N__26615\
        );

    \I__3440\ : CEMux
    port map (
            O => \N__26625\,
            I => \N__26615\
        );

    \I__3439\ : CEMux
    port map (
            O => \N__26624\,
            I => \N__26615\
        );

    \I__3438\ : GlobalMux
    port map (
            O => \N__26615\,
            I => \N__26612\
        );

    \I__3437\ : gio2CtrlBuf
    port map (
            O => \N__26612\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0_g\
        );

    \I__3436\ : IoInMux
    port map (
            O => \N__26609\,
            I => \N__26606\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__26606\,
            I => \N__26603\
        );

    \I__3434\ : Odrv12
    port map (
            O => \N__26603\,
            I => s4_phy_c
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__26600\,
            I => \N__26596\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__26599\,
            I => \N__26592\
        );

    \I__3431\ : InMux
    port map (
            O => \N__26596\,
            I => \N__26589\
        );

    \I__3430\ : InMux
    port map (
            O => \N__26595\,
            I => \N__26586\
        );

    \I__3429\ : InMux
    port map (
            O => \N__26592\,
            I => \N__26583\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__26589\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__26586\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__26583\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__3425\ : InMux
    port map (
            O => \N__26576\,
            I => \N__26572\
        );

    \I__3424\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26569\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__26572\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__26569\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__3421\ : InMux
    port map (
            O => \N__26564\,
            I => \N__26561\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__26561\,
            I => \phase_controller_inst2.state_ns_0_0_1\
        );

    \I__3419\ : InMux
    port map (
            O => \N__26558\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_19\
        );

    \I__3418\ : InMux
    port map (
            O => \N__26555\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_20\
        );

    \I__3417\ : InMux
    port map (
            O => \N__26552\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_21\
        );

    \I__3416\ : InMux
    port map (
            O => \N__26549\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_22\
        );

    \I__3415\ : InMux
    port map (
            O => \N__26546\,
            I => \bfn_8_23_0_\
        );

    \I__3414\ : InMux
    port map (
            O => \N__26543\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_24\
        );

    \I__3413\ : InMux
    port map (
            O => \N__26540\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_25\
        );

    \I__3412\ : InMux
    port map (
            O => \N__26537\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_26\
        );

    \I__3411\ : InMux
    port map (
            O => \N__26534\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_27\
        );

    \I__3410\ : InMux
    port map (
            O => \N__26531\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_10\
        );

    \I__3409\ : InMux
    port map (
            O => \N__26528\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_11\
        );

    \I__3408\ : InMux
    port map (
            O => \N__26525\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_12\
        );

    \I__3407\ : InMux
    port map (
            O => \N__26522\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_13\
        );

    \I__3406\ : InMux
    port map (
            O => \N__26519\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_14\
        );

    \I__3405\ : InMux
    port map (
            O => \N__26516\,
            I => \bfn_8_22_0_\
        );

    \I__3404\ : InMux
    port map (
            O => \N__26513\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_16\
        );

    \I__3403\ : CascadeMux
    port map (
            O => \N__26510\,
            I => \N__26506\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__26509\,
            I => \N__26503\
        );

    \I__3401\ : InMux
    port map (
            O => \N__26506\,
            I => \N__26497\
        );

    \I__3400\ : InMux
    port map (
            O => \N__26503\,
            I => \N__26497\
        );

    \I__3399\ : InMux
    port map (
            O => \N__26502\,
            I => \N__26494\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__26497\,
            I => \N__26491\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__26494\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_18\
        );

    \I__3396\ : Odrv4
    port map (
            O => \N__26491\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_18\
        );

    \I__3395\ : InMux
    port map (
            O => \N__26486\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_17\
        );

    \I__3394\ : InMux
    port map (
            O => \N__26483\,
            I => \N__26476\
        );

    \I__3393\ : InMux
    port map (
            O => \N__26482\,
            I => \N__26476\
        );

    \I__3392\ : InMux
    port map (
            O => \N__26481\,
            I => \N__26473\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__26476\,
            I => \N__26470\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__26473\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_19\
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__26470\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_19\
        );

    \I__3388\ : InMux
    port map (
            O => \N__26465\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_18\
        );

    \I__3387\ : InMux
    port map (
            O => \N__26462\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_1\
        );

    \I__3386\ : InMux
    port map (
            O => \N__26459\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_2\
        );

    \I__3385\ : InMux
    port map (
            O => \N__26456\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_3\
        );

    \I__3384\ : InMux
    port map (
            O => \N__26453\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_4\
        );

    \I__3383\ : InMux
    port map (
            O => \N__26450\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_5\
        );

    \I__3382\ : InMux
    port map (
            O => \N__26447\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_6\
        );

    \I__3381\ : InMux
    port map (
            O => \N__26444\,
            I => \bfn_8_21_0_\
        );

    \I__3380\ : InMux
    port map (
            O => \N__26441\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_8\
        );

    \I__3379\ : InMux
    port map (
            O => \N__26438\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_9\
        );

    \I__3378\ : InMux
    port map (
            O => \N__26435\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21\
        );

    \I__3377\ : InMux
    port map (
            O => \N__26432\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22\
        );

    \I__3376\ : InMux
    port map (
            O => \N__26429\,
            I => \bfn_8_19_0_\
        );

    \I__3375\ : InMux
    port map (
            O => \N__26426\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24\
        );

    \I__3374\ : InMux
    port map (
            O => \N__26423\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25\
        );

    \I__3373\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26417\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__26417\,
            I => \N__26413\
        );

    \I__3371\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26410\
        );

    \I__3370\ : Span4Mux_v
    port map (
            O => \N__26413\,
            I => \N__26405\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__26410\,
            I => \N__26405\
        );

    \I__3368\ : Odrv4
    port map (
            O => \N__26405\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_27
        );

    \I__3367\ : InMux
    port map (
            O => \N__26402\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26\
        );

    \I__3366\ : InMux
    port map (
            O => \N__26399\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27\
        );

    \I__3365\ : InMux
    port map (
            O => \N__26396\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_0\
        );

    \I__3364\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26390\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__26390\,
            I => \N__26387\
        );

    \I__3362\ : Span4Mux_h
    port map (
            O => \N__26387\,
            I => \N__26383\
        );

    \I__3361\ : InMux
    port map (
            O => \N__26386\,
            I => \N__26380\
        );

    \I__3360\ : Odrv4
    port map (
            O => \N__26383\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_13
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__26380\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_13
        );

    \I__3358\ : InMux
    port map (
            O => \N__26375\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12\
        );

    \I__3357\ : InMux
    port map (
            O => \N__26372\,
            I => \N__26369\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__26369\,
            I => \N__26366\
        );

    \I__3355\ : Span4Mux_h
    port map (
            O => \N__26366\,
            I => \N__26362\
        );

    \I__3354\ : InMux
    port map (
            O => \N__26365\,
            I => \N__26359\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__26362\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_14
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__26359\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_14
        );

    \I__3351\ : InMux
    port map (
            O => \N__26354\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13\
        );

    \I__3350\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26348\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__26348\,
            I => \N__26345\
        );

    \I__3348\ : Span4Mux_v
    port map (
            O => \N__26345\,
            I => \N__26341\
        );

    \I__3347\ : InMux
    port map (
            O => \N__26344\,
            I => \N__26338\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__26341\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_15
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__26338\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_15
        );

    \I__3344\ : InMux
    port map (
            O => \N__26333\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14\
        );

    \I__3343\ : InMux
    port map (
            O => \N__26330\,
            I => \N__26326\
        );

    \I__3342\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26323\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__26326\,
            I => \N__26320\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__26323\,
            I => \N__26317\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__26320\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_16
        );

    \I__3338\ : Odrv4
    port map (
            O => \N__26317\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_16
        );

    \I__3337\ : InMux
    port map (
            O => \N__26312\,
            I => \bfn_8_18_0_\
        );

    \I__3336\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26305\
        );

    \I__3335\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26302\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__26305\,
            I => \N__26299\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__26302\,
            I => \N__26296\
        );

    \I__3332\ : Odrv4
    port map (
            O => \N__26299\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_17
        );

    \I__3331\ : Odrv4
    port map (
            O => \N__26296\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_17
        );

    \I__3330\ : InMux
    port map (
            O => \N__26291\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16\
        );

    \I__3329\ : InMux
    port map (
            O => \N__26288\,
            I => \N__26285\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__26285\,
            I => \N__26281\
        );

    \I__3327\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26278\
        );

    \I__3326\ : Span4Mux_v
    port map (
            O => \N__26281\,
            I => \N__26273\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__26278\,
            I => \N__26273\
        );

    \I__3324\ : Odrv4
    port map (
            O => \N__26273\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_18
        );

    \I__3323\ : InMux
    port map (
            O => \N__26270\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17\
        );

    \I__3322\ : InMux
    port map (
            O => \N__26267\,
            I => \N__26264\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__26264\,
            I => \N__26260\
        );

    \I__3320\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26257\
        );

    \I__3319\ : Span4Mux_v
    port map (
            O => \N__26260\,
            I => \N__26252\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__26257\,
            I => \N__26252\
        );

    \I__3317\ : Odrv4
    port map (
            O => \N__26252\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_19
        );

    \I__3316\ : InMux
    port map (
            O => \N__26249\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18\
        );

    \I__3315\ : InMux
    port map (
            O => \N__26246\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19\
        );

    \I__3314\ : InMux
    port map (
            O => \N__26243\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20\
        );

    \I__3313\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26237\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__26237\,
            I => \N__26233\
        );

    \I__3311\ : InMux
    port map (
            O => \N__26236\,
            I => \N__26230\
        );

    \I__3310\ : Odrv4
    port map (
            O => \N__26233\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_5
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__26230\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_5
        );

    \I__3308\ : InMux
    port map (
            O => \N__26225\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4\
        );

    \I__3307\ : InMux
    port map (
            O => \N__26222\,
            I => \N__26219\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__26219\,
            I => \N__26215\
        );

    \I__3305\ : InMux
    port map (
            O => \N__26218\,
            I => \N__26212\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__26215\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_6
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__26212\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_6
        );

    \I__3302\ : InMux
    port map (
            O => \N__26207\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5\
        );

    \I__3301\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26200\
        );

    \I__3300\ : InMux
    port map (
            O => \N__26203\,
            I => \N__26197\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__26200\,
            I => \N__26194\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__26197\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_7
        );

    \I__3297\ : Odrv4
    port map (
            O => \N__26194\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_7
        );

    \I__3296\ : InMux
    port map (
            O => \N__26189\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6\
        );

    \I__3295\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26182\
        );

    \I__3294\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26179\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__26182\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_8
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__26179\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_8
        );

    \I__3291\ : InMux
    port map (
            O => \N__26174\,
            I => \bfn_8_17_0_\
        );

    \I__3290\ : InMux
    port map (
            O => \N__26171\,
            I => \N__26168\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__26168\,
            I => \N__26164\
        );

    \I__3288\ : InMux
    port map (
            O => \N__26167\,
            I => \N__26161\
        );

    \I__3287\ : Odrv4
    port map (
            O => \N__26164\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_9
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__26161\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_9
        );

    \I__3285\ : InMux
    port map (
            O => \N__26156\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8\
        );

    \I__3284\ : InMux
    port map (
            O => \N__26153\,
            I => \N__26149\
        );

    \I__3283\ : InMux
    port map (
            O => \N__26152\,
            I => \N__26146\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__26149\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_10
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__26146\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_10
        );

    \I__3280\ : InMux
    port map (
            O => \N__26141\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9\
        );

    \I__3279\ : InMux
    port map (
            O => \N__26138\,
            I => \N__26135\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__26135\,
            I => \N__26131\
        );

    \I__3277\ : InMux
    port map (
            O => \N__26134\,
            I => \N__26128\
        );

    \I__3276\ : Odrv4
    port map (
            O => \N__26131\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_11
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__26128\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_11
        );

    \I__3274\ : InMux
    port map (
            O => \N__26123\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10\
        );

    \I__3273\ : InMux
    port map (
            O => \N__26120\,
            I => \N__26117\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__26117\,
            I => \N__26114\
        );

    \I__3271\ : Span4Mux_h
    port map (
            O => \N__26114\,
            I => \N__26110\
        );

    \I__3270\ : InMux
    port map (
            O => \N__26113\,
            I => \N__26107\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__26110\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_12
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__26107\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_12
        );

    \I__3267\ : InMux
    port map (
            O => \N__26102\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11\
        );

    \I__3266\ : InMux
    port map (
            O => \N__26099\,
            I => \N__26096\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__26096\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__3264\ : CascadeMux
    port map (
            O => \N__26093\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\
        );

    \I__3263\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26086\
        );

    \I__3262\ : InMux
    port map (
            O => \N__26089\,
            I => \N__26083\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__26086\,
            I => \N__26080\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__26083\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__3259\ : Odrv4
    port map (
            O => \N__26080\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__26075\,
            I => \N__26072\
        );

    \I__3257\ : InMux
    port map (
            O => \N__26072\,
            I => \N__26069\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__26069\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt30\
        );

    \I__3255\ : InMux
    port map (
            O => \N__26066\,
            I => \N__26063\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__26063\,
            I => \phase_controller_inst1.stoper_tr.measured_delay_tr_i_31\
        );

    \I__3253\ : InMux
    port map (
            O => \N__26060\,
            I => \N__26056\
        );

    \I__3252\ : InMux
    port map (
            O => \N__26059\,
            I => \N__26053\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__26056\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_1
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__26053\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_1
        );

    \I__3249\ : InMux
    port map (
            O => \N__26048\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0\
        );

    \I__3248\ : InMux
    port map (
            O => \N__26045\,
            I => \N__26042\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__26042\,
            I => \N__26038\
        );

    \I__3246\ : InMux
    port map (
            O => \N__26041\,
            I => \N__26035\
        );

    \I__3245\ : Odrv4
    port map (
            O => \N__26038\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_2
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__26035\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_2
        );

    \I__3243\ : InMux
    port map (
            O => \N__26030\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1\
        );

    \I__3242\ : InMux
    port map (
            O => \N__26027\,
            I => \N__26023\
        );

    \I__3241\ : InMux
    port map (
            O => \N__26026\,
            I => \N__26020\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__26023\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_3
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__26020\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_3
        );

    \I__3238\ : InMux
    port map (
            O => \N__26015\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2\
        );

    \I__3237\ : InMux
    port map (
            O => \N__26012\,
            I => \N__26009\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__26009\,
            I => \N__26005\
        );

    \I__3235\ : InMux
    port map (
            O => \N__26008\,
            I => \N__26002\
        );

    \I__3234\ : Odrv4
    port map (
            O => \N__26005\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_4
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__26002\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_4
        );

    \I__3232\ : InMux
    port map (
            O => \N__25997\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3\
        );

    \I__3231\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25991\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25988\
        );

    \I__3229\ : Odrv4
    port map (
            O => \N__25988\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24\
        );

    \I__3228\ : CascadeMux
    port map (
            O => \N__25985\,
            I => \N__25982\
        );

    \I__3227\ : InMux
    port map (
            O => \N__25982\,
            I => \N__25979\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__25979\,
            I => \N__25976\
        );

    \I__3225\ : Span4Mux_h
    port map (
            O => \N__25976\,
            I => \N__25973\
        );

    \I__3224\ : Odrv4
    port map (
            O => \N__25973\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt24\
        );

    \I__3223\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25967\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__25967\,
            I => \N__25964\
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__25964\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt26\
        );

    \I__3220\ : CascadeMux
    port map (
            O => \N__25961\,
            I => \N__25958\
        );

    \I__3219\ : InMux
    port map (
            O => \N__25958\,
            I => \N__25955\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__25955\,
            I => \N__25952\
        );

    \I__3217\ : Span4Mux_v
    port map (
            O => \N__25952\,
            I => \N__25949\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__25949\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26\
        );

    \I__3215\ : InMux
    port map (
            O => \N__25946\,
            I => \bfn_8_15_0_\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__25943\,
            I => \N__25940\
        );

    \I__3213\ : InMux
    port map (
            O => \N__25940\,
            I => \N__25937\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__25937\,
            I => \N__25934\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__25934\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt28\
        );

    \I__3210\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25925\
        );

    \I__3209\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25925\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__25925\,
            I => \N__25921\
        );

    \I__3207\ : InMux
    port map (
            O => \N__25924\,
            I => \N__25918\
        );

    \I__3206\ : Span4Mux_v
    port map (
            O => \N__25921\,
            I => \N__25915\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__25918\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_29\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__25915\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_29\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__25910\,
            I => \N__25907\
        );

    \I__3202\ : InMux
    port map (
            O => \N__25907\,
            I => \N__25901\
        );

    \I__3201\ : InMux
    port map (
            O => \N__25906\,
            I => \N__25901\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__25901\,
            I => \N__25897\
        );

    \I__3199\ : InMux
    port map (
            O => \N__25900\,
            I => \N__25894\
        );

    \I__3198\ : Span4Mux_v
    port map (
            O => \N__25897\,
            I => \N__25891\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__25894\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_28\
        );

    \I__3196\ : Odrv4
    port map (
            O => \N__25891\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_28\
        );

    \I__3195\ : InMux
    port map (
            O => \N__25886\,
            I => \N__25883\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__25883\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28\
        );

    \I__3193\ : InMux
    port map (
            O => \N__25880\,
            I => \N__25877\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__25877\,
            I => \N__25870\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__25876\,
            I => \N__25867\
        );

    \I__3190\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25861\
        );

    \I__3189\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25861\
        );

    \I__3188\ : InMux
    port map (
            O => \N__25873\,
            I => \N__25858\
        );

    \I__3187\ : Span4Mux_v
    port map (
            O => \N__25870\,
            I => \N__25855\
        );

    \I__3186\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25852\
        );

    \I__3185\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25849\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__25861\,
            I => \N__25846\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__25858\,
            I => \N__25843\
        );

    \I__3182\ : Span4Mux_v
    port map (
            O => \N__25855\,
            I => \N__25840\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__25852\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__25849\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__25846\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__3178\ : Odrv4
    port map (
            O => \N__25843\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__25840\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__3176\ : InMux
    port map (
            O => \N__25829\,
            I => \N__25823\
        );

    \I__3175\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25823\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__25823\,
            I => \N__25820\
        );

    \I__3173\ : Span12Mux_s10_v
    port map (
            O => \N__25820\,
            I => \N__25816\
        );

    \I__3172\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25813\
        );

    \I__3171\ : Odrv12
    port map (
            O => \N__25816\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__25813\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__25808\,
            I => \N__25804\
        );

    \I__3168\ : InMux
    port map (
            O => \N__25807\,
            I => \N__25801\
        );

    \I__3167\ : InMux
    port map (
            O => \N__25804\,
            I => \N__25798\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__25801\,
            I => \N__25795\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__25798\,
            I => \N__25792\
        );

    \I__3164\ : Span4Mux_v
    port map (
            O => \N__25795\,
            I => \N__25787\
        );

    \I__3163\ : Span4Mux_v
    port map (
            O => \N__25792\,
            I => \N__25787\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__25787\,
            I => \phase_controller_inst2.stoper_tr.counter\
        );

    \I__3161\ : InMux
    port map (
            O => \N__25784\,
            I => \N__25781\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__25781\,
            I => \N__25778\
        );

    \I__3159\ : Span4Mux_h
    port map (
            O => \N__25778\,
            I => \N__25775\
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__25775\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_12\
        );

    \I__3157\ : InMux
    port map (
            O => \N__25772\,
            I => \N__25768\
        );

    \I__3156\ : InMux
    port map (
            O => \N__25771\,
            I => \N__25765\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__25768\,
            I => \N__25762\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__25765\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_12\
        );

    \I__3153\ : Odrv12
    port map (
            O => \N__25762\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_12\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__25757\,
            I => \N__25754\
        );

    \I__3151\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25751\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__25751\,
            I => \phase_controller_inst2.stoper_tr.counter_i_12\
        );

    \I__3149\ : InMux
    port map (
            O => \N__25748\,
            I => \N__25744\
        );

    \I__3148\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25741\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__25744\,
            I => \N__25738\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__25741\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_13\
        );

    \I__3145\ : Odrv12
    port map (
            O => \N__25738\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_13\
        );

    \I__3144\ : InMux
    port map (
            O => \N__25733\,
            I => \N__25730\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__25730\,
            I => \N__25727\
        );

    \I__3142\ : Span4Mux_v
    port map (
            O => \N__25727\,
            I => \N__25724\
        );

    \I__3141\ : Odrv4
    port map (
            O => \N__25724\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_13\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__25721\,
            I => \N__25718\
        );

    \I__3139\ : InMux
    port map (
            O => \N__25718\,
            I => \N__25715\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__25715\,
            I => \N__25712\
        );

    \I__3137\ : Odrv4
    port map (
            O => \N__25712\,
            I => \phase_controller_inst2.stoper_tr.counter_i_13\
        );

    \I__3136\ : InMux
    port map (
            O => \N__25709\,
            I => \N__25705\
        );

    \I__3135\ : InMux
    port map (
            O => \N__25708\,
            I => \N__25702\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__25705\,
            I => \N__25699\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__25702\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_14\
        );

    \I__3132\ : Odrv12
    port map (
            O => \N__25699\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_14\
        );

    \I__3131\ : InMux
    port map (
            O => \N__25694\,
            I => \N__25691\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__25691\,
            I => \N__25688\
        );

    \I__3129\ : Span4Mux_h
    port map (
            O => \N__25688\,
            I => \N__25685\
        );

    \I__3128\ : Odrv4
    port map (
            O => \N__25685\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_14\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__25682\,
            I => \N__25679\
        );

    \I__3126\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25676\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__25676\,
            I => \phase_controller_inst2.stoper_tr.counter_i_14\
        );

    \I__3124\ : InMux
    port map (
            O => \N__25673\,
            I => \N__25670\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__25670\,
            I => \N__25666\
        );

    \I__3122\ : InMux
    port map (
            O => \N__25669\,
            I => \N__25663\
        );

    \I__3121\ : Span4Mux_v
    port map (
            O => \N__25666\,
            I => \N__25660\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__25663\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_15\
        );

    \I__3119\ : Odrv4
    port map (
            O => \N__25660\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_15\
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__25655\,
            I => \N__25652\
        );

    \I__3117\ : InMux
    port map (
            O => \N__25652\,
            I => \N__25649\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__25649\,
            I => \N__25646\
        );

    \I__3115\ : Span4Mux_v
    port map (
            O => \N__25646\,
            I => \N__25643\
        );

    \I__3114\ : Odrv4
    port map (
            O => \N__25643\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_15\
        );

    \I__3113\ : InMux
    port map (
            O => \N__25640\,
            I => \N__25637\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__25637\,
            I => \phase_controller_inst2.stoper_tr.counter_i_15\
        );

    \I__3111\ : InMux
    port map (
            O => \N__25634\,
            I => \N__25631\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__25631\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt16\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__25628\,
            I => \N__25625\
        );

    \I__3108\ : InMux
    port map (
            O => \N__25625\,
            I => \N__25622\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__25622\,
            I => \N__25619\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__25619\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16\
        );

    \I__3105\ : InMux
    port map (
            O => \N__25616\,
            I => \N__25613\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__25613\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__25610\,
            I => \N__25607\
        );

    \I__3102\ : InMux
    port map (
            O => \N__25607\,
            I => \N__25604\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__25604\,
            I => \N__25601\
        );

    \I__3100\ : Odrv4
    port map (
            O => \N__25601\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt18\
        );

    \I__3099\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25595\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__25595\,
            I => \N__25592\
        );

    \I__3097\ : Span4Mux_h
    port map (
            O => \N__25592\,
            I => \N__25589\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__25589\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__25586\,
            I => \N__25583\
        );

    \I__3094\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25580\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__25580\,
            I => \N__25577\
        );

    \I__3092\ : Span4Mux_v
    port map (
            O => \N__25577\,
            I => \N__25574\
        );

    \I__3091\ : Odrv4
    port map (
            O => \N__25574\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt20\
        );

    \I__3090\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25568\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__25568\,
            I => \N__25565\
        );

    \I__3088\ : Odrv4
    port map (
            O => \N__25565\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__25562\,
            I => \N__25559\
        );

    \I__3086\ : InMux
    port map (
            O => \N__25559\,
            I => \N__25556\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__25556\,
            I => \N__25553\
        );

    \I__3084\ : Span4Mux_v
    port map (
            O => \N__25553\,
            I => \N__25550\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__25550\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt22\
        );

    \I__3082\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25543\
        );

    \I__3081\ : InMux
    port map (
            O => \N__25546\,
            I => \N__25540\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__25543\,
            I => \N__25537\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__25540\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_5\
        );

    \I__3078\ : Odrv12
    port map (
            O => \N__25537\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_5\
        );

    \I__3077\ : InMux
    port map (
            O => \N__25532\,
            I => \N__25529\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__25529\,
            I => \N__25526\
        );

    \I__3075\ : Span4Mux_h
    port map (
            O => \N__25526\,
            I => \N__25523\
        );

    \I__3074\ : Odrv4
    port map (
            O => \N__25523\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_5\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__25520\,
            I => \N__25517\
        );

    \I__3072\ : InMux
    port map (
            O => \N__25517\,
            I => \N__25514\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__25514\,
            I => \phase_controller_inst2.stoper_tr.counter_i_5\
        );

    \I__3070\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25508\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__25508\,
            I => \N__25505\
        );

    \I__3068\ : Span4Mux_v
    port map (
            O => \N__25505\,
            I => \N__25502\
        );

    \I__3067\ : Odrv4
    port map (
            O => \N__25502\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_6\
        );

    \I__3066\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25496\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__25496\,
            I => \N__25492\
        );

    \I__3064\ : InMux
    port map (
            O => \N__25495\,
            I => \N__25489\
        );

    \I__3063\ : Span4Mux_v
    port map (
            O => \N__25492\,
            I => \N__25486\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__25489\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_6\
        );

    \I__3061\ : Odrv4
    port map (
            O => \N__25486\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_6\
        );

    \I__3060\ : CascadeMux
    port map (
            O => \N__25481\,
            I => \N__25478\
        );

    \I__3059\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25475\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__25475\,
            I => \N__25472\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__25472\,
            I => \phase_controller_inst2.stoper_tr.counter_i_6\
        );

    \I__3056\ : InMux
    port map (
            O => \N__25469\,
            I => \N__25466\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__25466\,
            I => \N__25463\
        );

    \I__3054\ : Odrv4
    port map (
            O => \N__25463\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_7\
        );

    \I__3053\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25457\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__25457\,
            I => \N__25453\
        );

    \I__3051\ : InMux
    port map (
            O => \N__25456\,
            I => \N__25450\
        );

    \I__3050\ : Span4Mux_v
    port map (
            O => \N__25453\,
            I => \N__25447\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__25450\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_7\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__25447\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_7\
        );

    \I__3047\ : CascadeMux
    port map (
            O => \N__25442\,
            I => \N__25439\
        );

    \I__3046\ : InMux
    port map (
            O => \N__25439\,
            I => \N__25436\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__25436\,
            I => \phase_controller_inst2.stoper_tr.counter_i_7\
        );

    \I__3044\ : InMux
    port map (
            O => \N__25433\,
            I => \N__25429\
        );

    \I__3043\ : InMux
    port map (
            O => \N__25432\,
            I => \N__25426\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__25429\,
            I => \N__25423\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__25426\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_8\
        );

    \I__3040\ : Odrv12
    port map (
            O => \N__25423\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_8\
        );

    \I__3039\ : InMux
    port map (
            O => \N__25418\,
            I => \N__25415\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__25415\,
            I => \N__25412\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__25412\,
            I => \N__25409\
        );

    \I__3036\ : Odrv4
    port map (
            O => \N__25409\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_8\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__25406\,
            I => \N__25403\
        );

    \I__3034\ : InMux
    port map (
            O => \N__25403\,
            I => \N__25400\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__25400\,
            I => \phase_controller_inst2.stoper_tr.counter_i_8\
        );

    \I__3032\ : InMux
    port map (
            O => \N__25397\,
            I => \N__25394\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__25394\,
            I => \N__25391\
        );

    \I__3030\ : Span4Mux_v
    port map (
            O => \N__25391\,
            I => \N__25388\
        );

    \I__3029\ : Odrv4
    port map (
            O => \N__25388\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_9\
        );

    \I__3028\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25381\
        );

    \I__3027\ : InMux
    port map (
            O => \N__25384\,
            I => \N__25378\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__25381\,
            I => \N__25375\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__25378\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_9\
        );

    \I__3024\ : Odrv12
    port map (
            O => \N__25375\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_9\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__25370\,
            I => \N__25367\
        );

    \I__3022\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25364\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__25364\,
            I => \phase_controller_inst2.stoper_tr.counter_i_9\
        );

    \I__3020\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25358\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__25358\,
            I => \N__25355\
        );

    \I__3018\ : Span4Mux_h
    port map (
            O => \N__25355\,
            I => \N__25352\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__25352\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_10\
        );

    \I__3016\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25345\
        );

    \I__3015\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25342\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__25345\,
            I => \N__25339\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__25342\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_10\
        );

    \I__3012\ : Odrv12
    port map (
            O => \N__25339\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_10\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__25334\,
            I => \N__25331\
        );

    \I__3010\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25328\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__25328\,
            I => \phase_controller_inst2.stoper_tr.counter_i_10\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__25325\,
            I => \N__25322\
        );

    \I__3007\ : InMux
    port map (
            O => \N__25322\,
            I => \N__25319\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__25319\,
            I => \N__25316\
        );

    \I__3005\ : Odrv4
    port map (
            O => \N__25316\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_11\
        );

    \I__3004\ : InMux
    port map (
            O => \N__25313\,
            I => \N__25309\
        );

    \I__3003\ : InMux
    port map (
            O => \N__25312\,
            I => \N__25306\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__25309\,
            I => \N__25303\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__25306\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_11\
        );

    \I__3000\ : Odrv12
    port map (
            O => \N__25303\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_11\
        );

    \I__2999\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25295\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__25295\,
            I => \phase_controller_inst2.stoper_tr.counter_i_11\
        );

    \I__2997\ : InMux
    port map (
            O => \N__25292\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_28\
        );

    \I__2996\ : InMux
    port map (
            O => \N__25289\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_29\
        );

    \I__2995\ : InMux
    port map (
            O => \N__25286\,
            I => \N__25246\
        );

    \I__2994\ : InMux
    port map (
            O => \N__25285\,
            I => \N__25246\
        );

    \I__2993\ : InMux
    port map (
            O => \N__25284\,
            I => \N__25246\
        );

    \I__2992\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25246\
        );

    \I__2991\ : InMux
    port map (
            O => \N__25282\,
            I => \N__25237\
        );

    \I__2990\ : InMux
    port map (
            O => \N__25281\,
            I => \N__25237\
        );

    \I__2989\ : InMux
    port map (
            O => \N__25280\,
            I => \N__25237\
        );

    \I__2988\ : InMux
    port map (
            O => \N__25279\,
            I => \N__25237\
        );

    \I__2987\ : InMux
    port map (
            O => \N__25278\,
            I => \N__25228\
        );

    \I__2986\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25228\
        );

    \I__2985\ : InMux
    port map (
            O => \N__25276\,
            I => \N__25228\
        );

    \I__2984\ : InMux
    port map (
            O => \N__25275\,
            I => \N__25228\
        );

    \I__2983\ : InMux
    port map (
            O => \N__25274\,
            I => \N__25219\
        );

    \I__2982\ : InMux
    port map (
            O => \N__25273\,
            I => \N__25219\
        );

    \I__2981\ : InMux
    port map (
            O => \N__25272\,
            I => \N__25219\
        );

    \I__2980\ : InMux
    port map (
            O => \N__25271\,
            I => \N__25219\
        );

    \I__2979\ : InMux
    port map (
            O => \N__25270\,
            I => \N__25210\
        );

    \I__2978\ : InMux
    port map (
            O => \N__25269\,
            I => \N__25210\
        );

    \I__2977\ : InMux
    port map (
            O => \N__25268\,
            I => \N__25210\
        );

    \I__2976\ : InMux
    port map (
            O => \N__25267\,
            I => \N__25210\
        );

    \I__2975\ : InMux
    port map (
            O => \N__25266\,
            I => \N__25201\
        );

    \I__2974\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25201\
        );

    \I__2973\ : InMux
    port map (
            O => \N__25264\,
            I => \N__25201\
        );

    \I__2972\ : InMux
    port map (
            O => \N__25263\,
            I => \N__25201\
        );

    \I__2971\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25192\
        );

    \I__2970\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25192\
        );

    \I__2969\ : InMux
    port map (
            O => \N__25260\,
            I => \N__25192\
        );

    \I__2968\ : InMux
    port map (
            O => \N__25259\,
            I => \N__25192\
        );

    \I__2967\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25183\
        );

    \I__2966\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25183\
        );

    \I__2965\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25183\
        );

    \I__2964\ : InMux
    port map (
            O => \N__25255\,
            I => \N__25183\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__25246\,
            I => \N__25176\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__25237\,
            I => \N__25176\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__25228\,
            I => \N__25176\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__25219\,
            I => \phase_controller_inst2.stoper_tr.start_latched_i_0\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__25210\,
            I => \phase_controller_inst2.stoper_tr.start_latched_i_0\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__25201\,
            I => \phase_controller_inst2.stoper_tr.start_latched_i_0\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__25192\,
            I => \phase_controller_inst2.stoper_tr.start_latched_i_0\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__25183\,
            I => \phase_controller_inst2.stoper_tr.start_latched_i_0\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__25176\,
            I => \phase_controller_inst2.stoper_tr.start_latched_i_0\
        );

    \I__2954\ : InMux
    port map (
            O => \N__25163\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_30\
        );

    \I__2953\ : CEMux
    port map (
            O => \N__25160\,
            I => \N__25148\
        );

    \I__2952\ : CEMux
    port map (
            O => \N__25159\,
            I => \N__25148\
        );

    \I__2951\ : CEMux
    port map (
            O => \N__25158\,
            I => \N__25148\
        );

    \I__2950\ : CEMux
    port map (
            O => \N__25157\,
            I => \N__25148\
        );

    \I__2949\ : GlobalMux
    port map (
            O => \N__25148\,
            I => \N__25145\
        );

    \I__2948\ : gio2CtrlBuf
    port map (
            O => \N__25145\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0_g\
        );

    \I__2947\ : InMux
    port map (
            O => \N__25142\,
            I => \N__25139\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__25139\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_0\
        );

    \I__2945\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25132\
        );

    \I__2944\ : InMux
    port map (
            O => \N__25135\,
            I => \N__25129\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__25132\,
            I => \N__25126\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__25129\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_0\
        );

    \I__2941\ : Odrv12
    port map (
            O => \N__25126\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_0\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__25121\,
            I => \N__25118\
        );

    \I__2939\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25115\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__25115\,
            I => \phase_controller_inst2.stoper_tr.counter_i_0\
        );

    \I__2937\ : InMux
    port map (
            O => \N__25112\,
            I => \N__25109\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__25109\,
            I => \N__25106\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__25106\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_1\
        );

    \I__2934\ : InMux
    port map (
            O => \N__25103\,
            I => \N__25099\
        );

    \I__2933\ : InMux
    port map (
            O => \N__25102\,
            I => \N__25096\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__25099\,
            I => \N__25093\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__25096\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_1\
        );

    \I__2930\ : Odrv12
    port map (
            O => \N__25093\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_1\
        );

    \I__2929\ : CascadeMux
    port map (
            O => \N__25088\,
            I => \N__25085\
        );

    \I__2928\ : InMux
    port map (
            O => \N__25085\,
            I => \N__25082\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__25082\,
            I => \phase_controller_inst2.stoper_tr.counter_i_1\
        );

    \I__2926\ : InMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__2924\ : Span4Mux_h
    port map (
            O => \N__25073\,
            I => \N__25070\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__25070\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_2\
        );

    \I__2922\ : InMux
    port map (
            O => \N__25067\,
            I => \N__25063\
        );

    \I__2921\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25060\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__25063\,
            I => \N__25057\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__25060\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_2\
        );

    \I__2918\ : Odrv12
    port map (
            O => \N__25057\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_2\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__25052\,
            I => \N__25049\
        );

    \I__2916\ : InMux
    port map (
            O => \N__25049\,
            I => \N__25046\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__25046\,
            I => \N__25043\
        );

    \I__2914\ : Odrv4
    port map (
            O => \N__25043\,
            I => \phase_controller_inst2.stoper_tr.counter_i_2\
        );

    \I__2913\ : InMux
    port map (
            O => \N__25040\,
            I => \N__25037\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__25037\,
            I => \N__25034\
        );

    \I__2911\ : Span4Mux_h
    port map (
            O => \N__25034\,
            I => \N__25031\
        );

    \I__2910\ : Odrv4
    port map (
            O => \N__25031\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_3\
        );

    \I__2909\ : InMux
    port map (
            O => \N__25028\,
            I => \N__25024\
        );

    \I__2908\ : InMux
    port map (
            O => \N__25027\,
            I => \N__25021\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__25024\,
            I => \N__25018\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__25021\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_3\
        );

    \I__2905\ : Odrv12
    port map (
            O => \N__25018\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_3\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__25013\,
            I => \N__25010\
        );

    \I__2903\ : InMux
    port map (
            O => \N__25010\,
            I => \N__25007\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__25007\,
            I => \phase_controller_inst2.stoper_tr.counter_i_3\
        );

    \I__2901\ : InMux
    port map (
            O => \N__25004\,
            I => \N__25001\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__25001\,
            I => \N__24998\
        );

    \I__2899\ : Span4Mux_h
    port map (
            O => \N__24998\,
            I => \N__24995\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__24995\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_4\
        );

    \I__2897\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24989\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__24989\,
            I => \N__24985\
        );

    \I__2895\ : InMux
    port map (
            O => \N__24988\,
            I => \N__24982\
        );

    \I__2894\ : Span4Mux_v
    port map (
            O => \N__24985\,
            I => \N__24979\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__24982\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_4\
        );

    \I__2892\ : Odrv4
    port map (
            O => \N__24979\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_4\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__24974\,
            I => \N__24971\
        );

    \I__2890\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24968\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__24968\,
            I => \N__24965\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__24965\,
            I => \phase_controller_inst2.stoper_tr.counter_i_4\
        );

    \I__2887\ : InMux
    port map (
            O => \N__24962\,
            I => \N__24957\
        );

    \I__2886\ : InMux
    port map (
            O => \N__24961\,
            I => \N__24952\
        );

    \I__2885\ : InMux
    port map (
            O => \N__24960\,
            I => \N__24952\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__24957\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_21\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__24952\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_21\
        );

    \I__2882\ : InMux
    port map (
            O => \N__24947\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_20\
        );

    \I__2881\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24939\
        );

    \I__2880\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24934\
        );

    \I__2879\ : InMux
    port map (
            O => \N__24942\,
            I => \N__24934\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__24939\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_22\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__24934\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_22\
        );

    \I__2876\ : InMux
    port map (
            O => \N__24929\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_21\
        );

    \I__2875\ : InMux
    port map (
            O => \N__24926\,
            I => \N__24921\
        );

    \I__2874\ : InMux
    port map (
            O => \N__24925\,
            I => \N__24916\
        );

    \I__2873\ : InMux
    port map (
            O => \N__24924\,
            I => \N__24916\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__24921\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_23\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__24916\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_23\
        );

    \I__2870\ : InMux
    port map (
            O => \N__24911\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_22\
        );

    \I__2869\ : InMux
    port map (
            O => \N__24908\,
            I => \N__24903\
        );

    \I__2868\ : InMux
    port map (
            O => \N__24907\,
            I => \N__24898\
        );

    \I__2867\ : InMux
    port map (
            O => \N__24906\,
            I => \N__24898\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__24903\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_24\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__24898\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_24\
        );

    \I__2864\ : InMux
    port map (
            O => \N__24893\,
            I => \bfn_8_11_0_\
        );

    \I__2863\ : InMux
    port map (
            O => \N__24890\,
            I => \N__24885\
        );

    \I__2862\ : InMux
    port map (
            O => \N__24889\,
            I => \N__24880\
        );

    \I__2861\ : InMux
    port map (
            O => \N__24888\,
            I => \N__24880\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__24885\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_25\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__24880\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_25\
        );

    \I__2858\ : InMux
    port map (
            O => \N__24875\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_24\
        );

    \I__2857\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24867\
        );

    \I__2856\ : InMux
    port map (
            O => \N__24871\,
            I => \N__24862\
        );

    \I__2855\ : InMux
    port map (
            O => \N__24870\,
            I => \N__24862\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__24867\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_26\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__24862\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_26\
        );

    \I__2852\ : InMux
    port map (
            O => \N__24857\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_25\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__24854\,
            I => \N__24849\
        );

    \I__2850\ : CascadeMux
    port map (
            O => \N__24853\,
            I => \N__24846\
        );

    \I__2849\ : InMux
    port map (
            O => \N__24852\,
            I => \N__24843\
        );

    \I__2848\ : InMux
    port map (
            O => \N__24849\,
            I => \N__24838\
        );

    \I__2847\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24838\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__24843\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_27\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__24838\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_27\
        );

    \I__2844\ : InMux
    port map (
            O => \N__24833\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_26\
        );

    \I__2843\ : InMux
    port map (
            O => \N__24830\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_27\
        );

    \I__2842\ : InMux
    port map (
            O => \N__24827\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_11\
        );

    \I__2841\ : InMux
    port map (
            O => \N__24824\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_12\
        );

    \I__2840\ : InMux
    port map (
            O => \N__24821\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_13\
        );

    \I__2839\ : InMux
    port map (
            O => \N__24818\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_14\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__24815\,
            I => \N__24811\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__24814\,
            I => \N__24808\
        );

    \I__2836\ : InMux
    port map (
            O => \N__24811\,
            I => \N__24803\
        );

    \I__2835\ : InMux
    port map (
            O => \N__24808\,
            I => \N__24803\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__24803\,
            I => \N__24799\
        );

    \I__2833\ : InMux
    port map (
            O => \N__24802\,
            I => \N__24796\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__24799\,
            I => \N__24793\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__24796\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_16\
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__24793\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_16\
        );

    \I__2829\ : InMux
    port map (
            O => \N__24788\,
            I => \bfn_8_10_0_\
        );

    \I__2828\ : InMux
    port map (
            O => \N__24785\,
            I => \N__24779\
        );

    \I__2827\ : InMux
    port map (
            O => \N__24784\,
            I => \N__24779\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__24779\,
            I => \N__24775\
        );

    \I__2825\ : InMux
    port map (
            O => \N__24778\,
            I => \N__24772\
        );

    \I__2824\ : Span4Mux_v
    port map (
            O => \N__24775\,
            I => \N__24769\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__24772\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_17\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__24769\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_17\
        );

    \I__2821\ : InMux
    port map (
            O => \N__24764\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_16\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__24761\,
            I => \N__24757\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__24760\,
            I => \N__24754\
        );

    \I__2818\ : InMux
    port map (
            O => \N__24757\,
            I => \N__24749\
        );

    \I__2817\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24749\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__24749\,
            I => \N__24745\
        );

    \I__2815\ : InMux
    port map (
            O => \N__24748\,
            I => \N__24742\
        );

    \I__2814\ : Span4Mux_v
    port map (
            O => \N__24745\,
            I => \N__24739\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__24742\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_18\
        );

    \I__2812\ : Odrv4
    port map (
            O => \N__24739\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_18\
        );

    \I__2811\ : InMux
    port map (
            O => \N__24734\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_17\
        );

    \I__2810\ : InMux
    port map (
            O => \N__24731\,
            I => \N__24725\
        );

    \I__2809\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24725\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__24725\,
            I => \N__24721\
        );

    \I__2807\ : InMux
    port map (
            O => \N__24724\,
            I => \N__24718\
        );

    \I__2806\ : Span4Mux_v
    port map (
            O => \N__24721\,
            I => \N__24715\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__24718\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_19\
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__24715\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_19\
        );

    \I__2803\ : InMux
    port map (
            O => \N__24710\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_18\
        );

    \I__2802\ : InMux
    port map (
            O => \N__24707\,
            I => \N__24702\
        );

    \I__2801\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24697\
        );

    \I__2800\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24697\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__24702\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_20\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__24697\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_20\
        );

    \I__2797\ : InMux
    port map (
            O => \N__24692\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_19\
        );

    \I__2796\ : InMux
    port map (
            O => \N__24689\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_2\
        );

    \I__2795\ : InMux
    port map (
            O => \N__24686\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_3\
        );

    \I__2794\ : InMux
    port map (
            O => \N__24683\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_4\
        );

    \I__2793\ : InMux
    port map (
            O => \N__24680\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_5\
        );

    \I__2792\ : InMux
    port map (
            O => \N__24677\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_6\
        );

    \I__2791\ : InMux
    port map (
            O => \N__24674\,
            I => \bfn_8_9_0_\
        );

    \I__2790\ : InMux
    port map (
            O => \N__24671\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_8\
        );

    \I__2789\ : InMux
    port map (
            O => \N__24668\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_9\
        );

    \I__2788\ : InMux
    port map (
            O => \N__24665\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_10\
        );

    \I__2787\ : CascadeMux
    port map (
            O => \N__24662\,
            I => \N__24659\
        );

    \I__2786\ : InMux
    port map (
            O => \N__24659\,
            I => \N__24656\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__24656\,
            I => \phase_controller_inst2.stoper_tr.un4_start_0\
        );

    \I__2784\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24644\
        );

    \I__2783\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24644\
        );

    \I__2782\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24644\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__24644\,
            I => \phase_controller_inst2.stateZ0Z_4\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__24641\,
            I => \N__24636\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__24640\,
            I => \N__24633\
        );

    \I__2778\ : InMux
    port map (
            O => \N__24639\,
            I => \N__24626\
        );

    \I__2777\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24626\
        );

    \I__2776\ : InMux
    port map (
            O => \N__24633\,
            I => \N__24626\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__24626\,
            I => \phase_controller_inst2.start_flagZ0\
        );

    \I__2774\ : InMux
    port map (
            O => \N__24623\,
            I => \N__24616\
        );

    \I__2773\ : InMux
    port map (
            O => \N__24622\,
            I => \N__24612\
        );

    \I__2772\ : InMux
    port map (
            O => \N__24621\,
            I => \N__24607\
        );

    \I__2771\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24607\
        );

    \I__2770\ : InMux
    port map (
            O => \N__24619\,
            I => \N__24604\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__24616\,
            I => \N__24601\
        );

    \I__2768\ : InMux
    port map (
            O => \N__24615\,
            I => \N__24598\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__24612\,
            I => \N__24595\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__24607\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__24604\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__24601\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__24598\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__24595\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__2761\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24577\
        );

    \I__2760\ : InMux
    port map (
            O => \N__24583\,
            I => \N__24577\
        );

    \I__2759\ : InMux
    port map (
            O => \N__24582\,
            I => \N__24574\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__24577\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__24574\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__2756\ : InMux
    port map (
            O => \N__24569\,
            I => \N__24566\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__24566\,
            I => \phase_controller_inst2.start_timer_tr_0_sqmuxa\
        );

    \I__2754\ : InMux
    port map (
            O => \N__24563\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_0\
        );

    \I__2753\ : InMux
    port map (
            O => \N__24560\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_1\
        );

    \I__2752\ : InMux
    port map (
            O => \N__24557\,
            I => \N__24551\
        );

    \I__2751\ : InMux
    port map (
            O => \N__24556\,
            I => \N__24551\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__24551\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_18\
        );

    \I__2749\ : InMux
    port map (
            O => \N__24548\,
            I => \N__24542\
        );

    \I__2748\ : InMux
    port map (
            O => \N__24547\,
            I => \N__24542\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__24542\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_19\
        );

    \I__2746\ : IoInMux
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__24536\,
            I => \N__24533\
        );

    \I__2744\ : Span4Mux_s1_v
    port map (
            O => \N__24533\,
            I => \N__24530\
        );

    \I__2743\ : Span4Mux_h
    port map (
            O => \N__24530\,
            I => \N__24527\
        );

    \I__2742\ : Odrv4
    port map (
            O => \N__24527\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__2741\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24518\
        );

    \I__2740\ : InMux
    port map (
            O => \N__24523\,
            I => \N__24518\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__24518\,
            I => \N__24515\
        );

    \I__2738\ : Odrv12
    port map (
            O => \N__24515\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_24\
        );

    \I__2737\ : InMux
    port map (
            O => \N__24512\,
            I => \N__24506\
        );

    \I__2736\ : InMux
    port map (
            O => \N__24511\,
            I => \N__24506\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__24506\,
            I => \N__24503\
        );

    \I__2734\ : Span12Mux_v
    port map (
            O => \N__24503\,
            I => \N__24500\
        );

    \I__2733\ : Odrv12
    port map (
            O => \N__24500\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_20\
        );

    \I__2732\ : InMux
    port map (
            O => \N__24497\,
            I => \N__24491\
        );

    \I__2731\ : InMux
    port map (
            O => \N__24496\,
            I => \N__24491\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__24491\,
            I => \N__24488\
        );

    \I__2729\ : Odrv12
    port map (
            O => \N__24488\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__24485\,
            I => \N__24481\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__24484\,
            I => \N__24478\
        );

    \I__2726\ : InMux
    port map (
            O => \N__24481\,
            I => \N__24473\
        );

    \I__2725\ : InMux
    port map (
            O => \N__24478\,
            I => \N__24473\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__24473\,
            I => \N__24470\
        );

    \I__2723\ : Span4Mux_v
    port map (
            O => \N__24470\,
            I => \N__24467\
        );

    \I__2722\ : Span4Mux_v
    port map (
            O => \N__24467\,
            I => \N__24464\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__24464\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_22\
        );

    \I__2720\ : CEMux
    port map (
            O => \N__24461\,
            I => \N__24458\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__24458\,
            I => \N__24452\
        );

    \I__2718\ : CEMux
    port map (
            O => \N__24457\,
            I => \N__24449\
        );

    \I__2717\ : CEMux
    port map (
            O => \N__24456\,
            I => \N__24444\
        );

    \I__2716\ : CEMux
    port map (
            O => \N__24455\,
            I => \N__24440\
        );

    \I__2715\ : Span4Mux_v
    port map (
            O => \N__24452\,
            I => \N__24432\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__24449\,
            I => \N__24432\
        );

    \I__2713\ : CEMux
    port map (
            O => \N__24448\,
            I => \N__24429\
        );

    \I__2712\ : CEMux
    port map (
            O => \N__24447\,
            I => \N__24426\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__24444\,
            I => \N__24423\
        );

    \I__2710\ : CEMux
    port map (
            O => \N__24443\,
            I => \N__24420\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__24440\,
            I => \N__24417\
        );

    \I__2708\ : CEMux
    port map (
            O => \N__24439\,
            I => \N__24414\
        );

    \I__2707\ : CEMux
    port map (
            O => \N__24438\,
            I => \N__24411\
        );

    \I__2706\ : CEMux
    port map (
            O => \N__24437\,
            I => \N__24408\
        );

    \I__2705\ : Span4Mux_h
    port map (
            O => \N__24432\,
            I => \N__24401\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__24429\,
            I => \N__24401\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__24426\,
            I => \N__24398\
        );

    \I__2702\ : Span4Mux_h
    port map (
            O => \N__24423\,
            I => \N__24395\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__24420\,
            I => \N__24392\
        );

    \I__2700\ : Span4Mux_h
    port map (
            O => \N__24417\,
            I => \N__24387\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__24414\,
            I => \N__24387\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__24411\,
            I => \N__24382\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__24408\,
            I => \N__24382\
        );

    \I__2696\ : CEMux
    port map (
            O => \N__24407\,
            I => \N__24379\
        );

    \I__2695\ : CEMux
    port map (
            O => \N__24406\,
            I => \N__24376\
        );

    \I__2694\ : Span4Mux_v
    port map (
            O => \N__24401\,
            I => \N__24373\
        );

    \I__2693\ : Span4Mux_v
    port map (
            O => \N__24398\,
            I => \N__24370\
        );

    \I__2692\ : Span4Mux_h
    port map (
            O => \N__24395\,
            I => \N__24365\
        );

    \I__2691\ : Span4Mux_h
    port map (
            O => \N__24392\,
            I => \N__24365\
        );

    \I__2690\ : Span4Mux_v
    port map (
            O => \N__24387\,
            I => \N__24356\
        );

    \I__2689\ : Span4Mux_v
    port map (
            O => \N__24382\,
            I => \N__24356\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__24379\,
            I => \N__24356\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__24376\,
            I => \N__24356\
        );

    \I__2686\ : Span4Mux_h
    port map (
            O => \N__24373\,
            I => \N__24353\
        );

    \I__2685\ : Span4Mux_v
    port map (
            O => \N__24370\,
            I => \N__24350\
        );

    \I__2684\ : Span4Mux_v
    port map (
            O => \N__24365\,
            I => \N__24347\
        );

    \I__2683\ : Span4Mux_v
    port map (
            O => \N__24356\,
            I => \N__24344\
        );

    \I__2682\ : Odrv4
    port map (
            O => \N__24353\,
            I => \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__2681\ : Odrv4
    port map (
            O => \N__24350\,
            I => \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__24347\,
            I => \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__24344\,
            I => \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__2678\ : InMux
    port map (
            O => \N__24335\,
            I => \N__24329\
        );

    \I__2677\ : InMux
    port map (
            O => \N__24334\,
            I => \N__24329\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__24329\,
            I => \N__24326\
        );

    \I__2675\ : Odrv12
    port map (
            O => \N__24326\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__24323\,
            I => \N__24319\
        );

    \I__2673\ : CascadeMux
    port map (
            O => \N__24322\,
            I => \N__24316\
        );

    \I__2672\ : InMux
    port map (
            O => \N__24319\,
            I => \N__24311\
        );

    \I__2671\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24311\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__24311\,
            I => \N__24308\
        );

    \I__2669\ : Odrv12
    port map (
            O => \N__24308\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_21\
        );

    \I__2668\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24299\
        );

    \I__2667\ : InMux
    port map (
            O => \N__24304\,
            I => \N__24299\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__24299\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_19\
        );

    \I__2665\ : InMux
    port map (
            O => \N__24296\,
            I => \N__24290\
        );

    \I__2664\ : InMux
    port map (
            O => \N__24295\,
            I => \N__24290\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__24290\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_18\
        );

    \I__2662\ : InMux
    port map (
            O => \N__24287\,
            I => \N__24281\
        );

    \I__2661\ : InMux
    port map (
            O => \N__24286\,
            I => \N__24281\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__24281\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_16\
        );

    \I__2659\ : InMux
    port map (
            O => \N__24278\,
            I => \N__24272\
        );

    \I__2658\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24272\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__24272\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_17\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__24269\,
            I => \N__24265\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__24268\,
            I => \N__24262\
        );

    \I__2654\ : InMux
    port map (
            O => \N__24265\,
            I => \N__24257\
        );

    \I__2653\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24257\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__24257\,
            I => \N__24254\
        );

    \I__2651\ : Span4Mux_h
    port map (
            O => \N__24254\,
            I => \N__24251\
        );

    \I__2650\ : Span4Mux_v
    port map (
            O => \N__24251\,
            I => \N__24248\
        );

    \I__2649\ : Odrv4
    port map (
            O => \N__24248\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_25\
        );

    \I__2648\ : CascadeMux
    port map (
            O => \N__24245\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31_cascade_\
        );

    \I__2647\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24239\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__24239\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__24236\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\
        );

    \I__2644\ : InMux
    port map (
            O => \N__24233\,
            I => \N__24227\
        );

    \I__2643\ : InMux
    port map (
            O => \N__24232\,
            I => \N__24227\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__24227\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_23\
        );

    \I__2641\ : InMux
    port map (
            O => \N__24224\,
            I => \N__24219\
        );

    \I__2640\ : InMux
    port map (
            O => \N__24223\,
            I => \N__24216\
        );

    \I__2639\ : InMux
    port map (
            O => \N__24222\,
            I => \N__24213\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__24219\,
            I => \N__24210\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__24216\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__24213\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__24210\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__24203\,
            I => \N__24200\
        );

    \I__2633\ : InMux
    port map (
            O => \N__24200\,
            I => \N__24197\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__24197\,
            I => \N__24194\
        );

    \I__2631\ : Odrv4
    port map (
            O => \N__24194\,
            I => \pwm_generator_inst.N_184_i\
        );

    \I__2630\ : InMux
    port map (
            O => \N__24191\,
            I => \N__24188\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__24188\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2628\ : InMux
    port map (
            O => \N__24185\,
            I => \N__24180\
        );

    \I__2627\ : InMux
    port map (
            O => \N__24184\,
            I => \N__24177\
        );

    \I__2626\ : InMux
    port map (
            O => \N__24183\,
            I => \N__24174\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__24180\,
            I => \N__24171\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__24177\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__24174\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__24171\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__24164\,
            I => \N__24161\
        );

    \I__2620\ : InMux
    port map (
            O => \N__24161\,
            I => \N__24158\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__24158\,
            I => \N__24155\
        );

    \I__2618\ : Span4Mux_h
    port map (
            O => \N__24155\,
            I => \N__24152\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__24152\,
            I => \pwm_generator_inst.N_185_i\
        );

    \I__2616\ : InMux
    port map (
            O => \N__24149\,
            I => \N__24146\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__24146\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2614\ : CascadeMux
    port map (
            O => \N__24143\,
            I => \N__24140\
        );

    \I__2613\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24137\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__24137\,
            I => \N__24134\
        );

    \I__2611\ : Span4Mux_v
    port map (
            O => \N__24134\,
            I => \N__24131\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__24131\,
            I => \pwm_generator_inst.N_186_i\
        );

    \I__2609\ : InMux
    port map (
            O => \N__24128\,
            I => \N__24123\
        );

    \I__2608\ : InMux
    port map (
            O => \N__24127\,
            I => \N__24120\
        );

    \I__2607\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24117\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__24123\,
            I => \N__24114\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__24120\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__24117\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__24114\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2602\ : InMux
    port map (
            O => \N__24107\,
            I => \N__24104\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__24104\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__24101\,
            I => \N__24098\
        );

    \I__2599\ : InMux
    port map (
            O => \N__24098\,
            I => \N__24095\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__24095\,
            I => \pwm_generator_inst.N_187_i\
        );

    \I__2597\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24088\
        );

    \I__2596\ : InMux
    port map (
            O => \N__24091\,
            I => \N__24084\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__24088\,
            I => \N__24081\
        );

    \I__2594\ : InMux
    port map (
            O => \N__24087\,
            I => \N__24078\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__24084\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2592\ : Odrv12
    port map (
            O => \N__24081\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__24078\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2590\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24068\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__24068\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__24065\,
            I => \N__24062\
        );

    \I__2587\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24059\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__24059\,
            I => \N__24056\
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__24056\,
            I => \pwm_generator_inst.N_188_i\
        );

    \I__2584\ : InMux
    port map (
            O => \N__24053\,
            I => \N__24049\
        );

    \I__2583\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24045\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__24049\,
            I => \N__24042\
        );

    \I__2581\ : InMux
    port map (
            O => \N__24048\,
            I => \N__24039\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__24045\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2579\ : Odrv12
    port map (
            O => \N__24042\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__24039\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2577\ : InMux
    port map (
            O => \N__24032\,
            I => \N__24029\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__24029\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2575\ : InMux
    port map (
            O => \N__24026\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2574\ : IoInMux
    port map (
            O => \N__24023\,
            I => \N__24020\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__24020\,
            I => \N__24017\
        );

    \I__2572\ : Span4Mux_s3_v
    port map (
            O => \N__24017\,
            I => \N__24014\
        );

    \I__2571\ : Sp12to4
    port map (
            O => \N__24014\,
            I => \N__24011\
        );

    \I__2570\ : Span12Mux_h
    port map (
            O => \N__24011\,
            I => \N__24008\
        );

    \I__2569\ : Span12Mux_v
    port map (
            O => \N__24008\,
            I => \N__24005\
        );

    \I__2568\ : Odrv12
    port map (
            O => \N__24005\,
            I => pwm_output_c
        );

    \I__2567\ : InMux
    port map (
            O => \N__24002\,
            I => \N__23999\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__23999\,
            I => \N__23995\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__23998\,
            I => \N__23992\
        );

    \I__2564\ : Span4Mux_h
    port map (
            O => \N__23995\,
            I => \N__23989\
        );

    \I__2563\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23986\
        );

    \I__2562\ : Odrv4
    port map (
            O => \N__23989\,
            I => \pwm_generator_inst.un18_threshold1_20\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__23986\,
            I => \pwm_generator_inst.un18_threshold1_20\
        );

    \I__2560\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23978\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__23978\,
            I => \pwm_generator_inst.un22_threshold_1_cry_2_THRU_CO\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__23975\,
            I => \N__23972\
        );

    \I__2557\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23969\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__23969\,
            I => \N__23966\
        );

    \I__2555\ : Span4Mux_v
    port map (
            O => \N__23966\,
            I => \N__23962\
        );

    \I__2554\ : InMux
    port map (
            O => \N__23965\,
            I => \N__23959\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__23962\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__23959\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0\
        );

    \I__2551\ : InMux
    port map (
            O => \N__23954\,
            I => \N__23951\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__23951\,
            I => \pwm_generator_inst.un22_threshold_1_cry_3_THRU_CO\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__23948\,
            I => \N__23945\
        );

    \I__2548\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23942\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__23942\,
            I => \N__23939\
        );

    \I__2546\ : Span4Mux_h
    port map (
            O => \N__23939\,
            I => \N__23935\
        );

    \I__2545\ : InMux
    port map (
            O => \N__23938\,
            I => \N__23932\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__23935\,
            I => \pwm_generator_inst.un18_threshold1_21\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__23932\,
            I => \pwm_generator_inst.un18_threshold1_21\
        );

    \I__2542\ : InMux
    port map (
            O => \N__23927\,
            I => \N__23924\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__23924\,
            I => \N__23921\
        );

    \I__2540\ : Span4Mux_h
    port map (
            O => \N__23921\,
            I => \N__23917\
        );

    \I__2539\ : InMux
    port map (
            O => \N__23920\,
            I => \N__23914\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__23917\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__23914\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0\
        );

    \I__2536\ : InMux
    port map (
            O => \N__23909\,
            I => \N__23906\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__23906\,
            I => \pwm_generator_inst.un22_threshold_1_cry_4_THRU_CO\
        );

    \I__2534\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23890\
        );

    \I__2533\ : InMux
    port map (
            O => \N__23902\,
            I => \N__23890\
        );

    \I__2532\ : InMux
    port map (
            O => \N__23901\,
            I => \N__23890\
        );

    \I__2531\ : InMux
    port map (
            O => \N__23900\,
            I => \N__23890\
        );

    \I__2530\ : CascadeMux
    port map (
            O => \N__23899\,
            I => \N__23886\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__23890\,
            I => \N__23881\
        );

    \I__2528\ : InMux
    port map (
            O => \N__23889\,
            I => \N__23876\
        );

    \I__2527\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23873\
        );

    \I__2526\ : InMux
    port map (
            O => \N__23885\,
            I => \N__23868\
        );

    \I__2525\ : InMux
    port map (
            O => \N__23884\,
            I => \N__23868\
        );

    \I__2524\ : Span4Mux_v
    port map (
            O => \N__23881\,
            I => \N__23865\
        );

    \I__2523\ : InMux
    port map (
            O => \N__23880\,
            I => \N__23860\
        );

    \I__2522\ : InMux
    port map (
            O => \N__23879\,
            I => \N__23860\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__23876\,
            I => \N__23857\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__23873\,
            I => \N__23852\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__23868\,
            I => \N__23852\
        );

    \I__2518\ : Span4Mux_v
    port map (
            O => \N__23865\,
            I => \N__23849\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__23860\,
            I => \N__23844\
        );

    \I__2516\ : Span4Mux_v
    port map (
            O => \N__23857\,
            I => \N__23844\
        );

    \I__2515\ : Odrv4
    port map (
            O => \N__23852\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1\
        );

    \I__2514\ : Odrv4
    port map (
            O => \N__23849\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__23844\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__23837\,
            I => \N__23834\
        );

    \I__2511\ : InMux
    port map (
            O => \N__23834\,
            I => \N__23831\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__23831\,
            I => \N__23827\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__23830\,
            I => \N__23824\
        );

    \I__2508\ : Span4Mux_h
    port map (
            O => \N__23827\,
            I => \N__23821\
        );

    \I__2507\ : InMux
    port map (
            O => \N__23824\,
            I => \N__23818\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__23821\,
            I => \pwm_generator_inst.un18_threshold1_22\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__23818\,
            I => \pwm_generator_inst.un18_threshold1_22\
        );

    \I__2504\ : InMux
    port map (
            O => \N__23813\,
            I => \N__23810\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__23810\,
            I => \N__23807\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__23807\,
            I => \N__23803\
        );

    \I__2501\ : InMux
    port map (
            O => \N__23806\,
            I => \N__23800\
        );

    \I__2500\ : Odrv4
    port map (
            O => \N__23803\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__23800\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__23795\,
            I => \N__23792\
        );

    \I__2497\ : InMux
    port map (
            O => \N__23792\,
            I => \N__23789\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__23789\,
            I => \pwm_generator_inst.N_179_i\
        );

    \I__2495\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23782\
        );

    \I__2494\ : InMux
    port map (
            O => \N__23785\,
            I => \N__23778\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__23782\,
            I => \N__23775\
        );

    \I__2492\ : InMux
    port map (
            O => \N__23781\,
            I => \N__23772\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__23778\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2490\ : Odrv12
    port map (
            O => \N__23775\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__23772\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2488\ : InMux
    port map (
            O => \N__23765\,
            I => \N__23762\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__23762\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2486\ : InMux
    port map (
            O => \N__23759\,
            I => \N__23755\
        );

    \I__2485\ : InMux
    port map (
            O => \N__23758\,
            I => \N__23751\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__23755\,
            I => \N__23748\
        );

    \I__2483\ : InMux
    port map (
            O => \N__23754\,
            I => \N__23745\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__23751\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2481\ : Odrv12
    port map (
            O => \N__23748\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__23745\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2479\ : CascadeMux
    port map (
            O => \N__23738\,
            I => \N__23735\
        );

    \I__2478\ : InMux
    port map (
            O => \N__23735\,
            I => \N__23732\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__23732\,
            I => \N__23729\
        );

    \I__2476\ : Span4Mux_h
    port map (
            O => \N__23729\,
            I => \N__23726\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__23726\,
            I => \pwm_generator_inst.N_180_i\
        );

    \I__2474\ : InMux
    port map (
            O => \N__23723\,
            I => \N__23720\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__23720\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__23717\,
            I => \N__23714\
        );

    \I__2471\ : InMux
    port map (
            O => \N__23714\,
            I => \N__23711\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__23711\,
            I => \pwm_generator_inst.N_181_i\
        );

    \I__2469\ : CascadeMux
    port map (
            O => \N__23708\,
            I => \N__23703\
        );

    \I__2468\ : InMux
    port map (
            O => \N__23707\,
            I => \N__23700\
        );

    \I__2467\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23697\
        );

    \I__2466\ : InMux
    port map (
            O => \N__23703\,
            I => \N__23694\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__23700\,
            I => \N__23691\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__23697\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__23694\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__23691\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2461\ : InMux
    port map (
            O => \N__23684\,
            I => \N__23681\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__23681\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2459\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23673\
        );

    \I__2458\ : InMux
    port map (
            O => \N__23677\,
            I => \N__23670\
        );

    \I__2457\ : InMux
    port map (
            O => \N__23676\,
            I => \N__23667\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__23673\,
            I => \N__23664\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__23670\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__23667\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__23664\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__23657\,
            I => \N__23654\
        );

    \I__2451\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23651\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__23651\,
            I => \pwm_generator_inst.N_182_i\
        );

    \I__2449\ : InMux
    port map (
            O => \N__23648\,
            I => \N__23645\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__23645\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__23642\,
            I => \N__23639\
        );

    \I__2446\ : InMux
    port map (
            O => \N__23639\,
            I => \N__23636\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__23636\,
            I => \pwm_generator_inst.N_183_i\
        );

    \I__2444\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23628\
        );

    \I__2443\ : InMux
    port map (
            O => \N__23632\,
            I => \N__23625\
        );

    \I__2442\ : InMux
    port map (
            O => \N__23631\,
            I => \N__23622\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__23628\,
            I => \N__23619\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__23625\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__23622\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2438\ : Odrv4
    port map (
            O => \N__23619\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2437\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__23609\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2435\ : InMux
    port map (
            O => \N__23606\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__2434\ : InMux
    port map (
            O => \N__23603\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__2433\ : InMux
    port map (
            O => \N__23600\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__2432\ : InMux
    port map (
            O => \N__23597\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__2431\ : InMux
    port map (
            O => \N__23594\,
            I => \bfn_3_13_0_\
        );

    \I__2430\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23573\
        );

    \I__2429\ : InMux
    port map (
            O => \N__23590\,
            I => \N__23573\
        );

    \I__2428\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23573\
        );

    \I__2427\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23573\
        );

    \I__2426\ : InMux
    port map (
            O => \N__23587\,
            I => \N__23568\
        );

    \I__2425\ : InMux
    port map (
            O => \N__23586\,
            I => \N__23568\
        );

    \I__2424\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23559\
        );

    \I__2423\ : InMux
    port map (
            O => \N__23584\,
            I => \N__23559\
        );

    \I__2422\ : InMux
    port map (
            O => \N__23583\,
            I => \N__23559\
        );

    \I__2421\ : InMux
    port map (
            O => \N__23582\,
            I => \N__23559\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__23573\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__23568\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__23559\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2417\ : InMux
    port map (
            O => \N__23552\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__2416\ : InMux
    port map (
            O => \N__23549\,
            I => \N__23546\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__23546\,
            I => \pwm_generator_inst.un22_threshold_1_cry_1_THRU_CO\
        );

    \I__2414\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23540\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__23540\,
            I => \N__23537\
        );

    \I__2412\ : Span4Mux_h
    port map (
            O => \N__23537\,
            I => \N__23533\
        );

    \I__2411\ : InMux
    port map (
            O => \N__23536\,
            I => \N__23530\
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__23533\,
            I => \pwm_generator_inst.un18_threshold1_19\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__23530\,
            I => \pwm_generator_inst.un18_threshold1_19\
        );

    \I__2408\ : CascadeMux
    port map (
            O => \N__23525\,
            I => \N__23522\
        );

    \I__2407\ : InMux
    port map (
            O => \N__23522\,
            I => \N__23516\
        );

    \I__2406\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23516\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__23516\,
            I => \N__23513\
        );

    \I__2404\ : Span4Mux_v
    port map (
            O => \N__23513\,
            I => \N__23510\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__23510\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRROZ0\
        );

    \I__2402\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23504\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__23504\,
            I => \N__23501\
        );

    \I__2400\ : Span4Mux_s3_h
    port map (
            O => \N__23501\,
            I => \N__23498\
        );

    \I__2399\ : Odrv4
    port map (
            O => \N__23498\,
            I => \pwm_generator_inst.un18_threshold_1_axb_19\
        );

    \I__2398\ : InMux
    port map (
            O => \N__23495\,
            I => \N__23489\
        );

    \I__2397\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23486\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__23493\,
            I => \N__23482\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__23492\,
            I => \N__23478\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__23489\,
            I => \N__23474\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__23486\,
            I => \N__23471\
        );

    \I__2392\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23460\
        );

    \I__2391\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23460\
        );

    \I__2390\ : InMux
    port map (
            O => \N__23481\,
            I => \N__23460\
        );

    \I__2389\ : InMux
    port map (
            O => \N__23478\,
            I => \N__23460\
        );

    \I__2388\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23460\
        );

    \I__2387\ : Span4Mux_h
    port map (
            O => \N__23474\,
            I => \N__23457\
        );

    \I__2386\ : Span12Mux_h
    port map (
            O => \N__23471\,
            I => \N__23454\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__23460\,
            I => \N__23451\
        );

    \I__2384\ : Span4Mux_v
    port map (
            O => \N__23457\,
            I => \N__23448\
        );

    \I__2383\ : Span12Mux_v
    port map (
            O => \N__23454\,
            I => \N__23445\
        );

    \I__2382\ : Span12Mux_h
    port map (
            O => \N__23451\,
            I => \N__23442\
        );

    \I__2381\ : Span4Mux_v
    port map (
            O => \N__23448\,
            I => \N__23439\
        );

    \I__2380\ : Odrv12
    port map (
            O => \N__23445\,
            I => \pwm_generator_inst.un5_threshold_1_26\
        );

    \I__2379\ : Odrv12
    port map (
            O => \N__23442\,
            I => \pwm_generator_inst.un5_threshold_1_26\
        );

    \I__2378\ : Odrv4
    port map (
            O => \N__23439\,
            I => \pwm_generator_inst.un5_threshold_1_26\
        );

    \I__2377\ : InMux
    port map (
            O => \N__23432\,
            I => \N__23429\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__23429\,
            I => \N__23426\
        );

    \I__2375\ : Span4Mux_h
    port map (
            O => \N__23426\,
            I => \N__23423\
        );

    \I__2374\ : Span4Mux_v
    port map (
            O => \N__23423\,
            I => \N__23420\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__23420\,
            I => \pwm_generator_inst.un5_threshold_2_1_16\
        );

    \I__2372\ : InMux
    port map (
            O => \N__23417\,
            I => \N__23414\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__23414\,
            I => \N__23411\
        );

    \I__2370\ : Span4Mux_v
    port map (
            O => \N__23411\,
            I => \N__23408\
        );

    \I__2369\ : Odrv4
    port map (
            O => \N__23408\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSONZ0\
        );

    \I__2368\ : InMux
    port map (
            O => \N__23405\,
            I => \N__23402\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__23402\,
            I => \N__23399\
        );

    \I__2366\ : Span4Mux_v
    port map (
            O => \N__23399\,
            I => \N__23395\
        );

    \I__2365\ : InMux
    port map (
            O => \N__23398\,
            I => \N__23392\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__23395\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__23392\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__23387\,
            I => \pwm_generator_inst.un5_threshold_add_1_axb_16Z0Z_1_cascade_\
        );

    \I__2361\ : InMux
    port map (
            O => \N__23384\,
            I => \N__23381\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__23381\,
            I => \N__23377\
        );

    \I__2359\ : InMux
    port map (
            O => \N__23380\,
            I => \N__23374\
        );

    \I__2358\ : Span4Mux_v
    port map (
            O => \N__23377\,
            I => \N__23371\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__23374\,
            I => \N__23368\
        );

    \I__2356\ : Span4Mux_v
    port map (
            O => \N__23371\,
            I => \N__23365\
        );

    \I__2355\ : Span4Mux_h
    port map (
            O => \N__23368\,
            I => \N__23362\
        );

    \I__2354\ : Odrv4
    port map (
            O => \N__23365\,
            I => \pwm_generator_inst.un5_threshold_2_1_15\
        );

    \I__2353\ : Odrv4
    port map (
            O => \N__23362\,
            I => \pwm_generator_inst.un5_threshold_2_1_15\
        );

    \I__2352\ : InMux
    port map (
            O => \N__23357\,
            I => \N__23354\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__23354\,
            I => \N__23351\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__23351\,
            I => \pwm_generator_inst.un5_threshold_add_1_axb_16\
        );

    \I__2349\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23345\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__23345\,
            I => \N__23341\
        );

    \I__2347\ : InMux
    port map (
            O => \N__23344\,
            I => \N__23338\
        );

    \I__2346\ : Odrv4
    port map (
            O => \N__23341\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__23338\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0\
        );

    \I__2344\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23330\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__23330\,
            I => \pwm_generator_inst.un18_threshold_1_axb_25\
        );

    \I__2342\ : InMux
    port map (
            O => \N__23327\,
            I => \N__23324\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__23324\,
            I => \N__23321\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__23321\,
            I => un8_start_stop
        );

    \I__2339\ : InMux
    port map (
            O => \N__23318\,
            I => \N__23315\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__2337\ : Glb2LocalMux
    port map (
            O => \N__23312\,
            I => \N__23309\
        );

    \I__2336\ : GlobalMux
    port map (
            O => \N__23309\,
            I => clk_12mhz
        );

    \I__2335\ : IoInMux
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__23303\,
            I => \N__23300\
        );

    \I__2333\ : Span4Mux_s0_v
    port map (
            O => \N__23300\,
            I => \N__23297\
        );

    \I__2332\ : Span4Mux_h
    port map (
            O => \N__23297\,
            I => \N__23294\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__23294\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__2330\ : InMux
    port map (
            O => \N__23291\,
            I => \bfn_3_12_0_\
        );

    \I__2329\ : InMux
    port map (
            O => \N__23288\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__2328\ : InMux
    port map (
            O => \N__23285\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__2327\ : InMux
    port map (
            O => \N__23282\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__2326\ : InMux
    port map (
            O => \N__23279\,
            I => \bfn_2_16_0_\
        );

    \I__2325\ : InMux
    port map (
            O => \N__23276\,
            I => \pwm_generator_inst.un22_threshold_1_cry_8\
        );

    \I__2324\ : InMux
    port map (
            O => \N__23273\,
            I => \N__23270\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__23270\,
            I => \pwm_generator_inst.un22_threshold_1_cry_8_THRU_CO\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__23267\,
            I => \N__23264\
        );

    \I__2321\ : InMux
    port map (
            O => \N__23264\,
            I => \N__23260\
        );

    \I__2320\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23257\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__23260\,
            I => \pwm_generator_inst.un18_threshold1_25\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__23257\,
            I => \pwm_generator_inst.un18_threshold1_25\
        );

    \I__2317\ : InMux
    port map (
            O => \N__23252\,
            I => \N__23249\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__23249\,
            I => \pwm_generator_inst.un22_threshold_1_cry_7_THRU_CO\
        );

    \I__2315\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23242\
        );

    \I__2314\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23239\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__23242\,
            I => \pwm_generator_inst.un22_threshold_1\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__23239\,
            I => \pwm_generator_inst.un22_threshold_1\
        );

    \I__2311\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23230\
        );

    \I__2310\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23227\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__23230\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__23227\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0\
        );

    \I__2307\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23219\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__23219\,
            I => \N__23216\
        );

    \I__2305\ : Odrv4
    port map (
            O => \N__23216\,
            I => \pwm_generator_inst.un22_threshold_1_cry_5_THRU_CO\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__23213\,
            I => \N__23210\
        );

    \I__2303\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23207\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__23207\,
            I => \N__23203\
        );

    \I__2301\ : InMux
    port map (
            O => \N__23206\,
            I => \N__23200\
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__23203\,
            I => \pwm_generator_inst.un18_threshold1_23\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__23200\,
            I => \pwm_generator_inst.un18_threshold1_23\
        );

    \I__2298\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23189\
        );

    \I__2297\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23189\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__23189\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0\
        );

    \I__2295\ : InMux
    port map (
            O => \N__23186\,
            I => \N__23183\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__23183\,
            I => \N__23180\
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__23180\,
            I => \pwm_generator_inst.un18_threshold_1_axb_23\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__23177\,
            I => \N__23173\
        );

    \I__2291\ : InMux
    port map (
            O => \N__23176\,
            I => \N__23170\
        );

    \I__2290\ : InMux
    port map (
            O => \N__23173\,
            I => \N__23167\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__23170\,
            I => \pwm_generator_inst.un18_threshold1_24\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__23167\,
            I => \pwm_generator_inst.un18_threshold1_24\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__23162\,
            I => \N__23159\
        );

    \I__2286\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23156\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__23156\,
            I => \N__23153\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__23153\,
            I => \pwm_generator_inst.un22_threshold_1_cry_6_THRU_CO\
        );

    \I__2283\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23144\
        );

    \I__2282\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23144\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__23144\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0\
        );

    \I__2280\ : InMux
    port map (
            O => \N__23141\,
            I => \N__23138\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__23138\,
            I => \pwm_generator_inst.un18_threshold_1_axb_24\
        );

    \I__2278\ : InMux
    port map (
            O => \N__23135\,
            I => \N__23132\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__23132\,
            I => \pwm_generator_inst.un1_counterlto2_0\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__23129\,
            I => \N__23126\
        );

    \I__2275\ : InMux
    port map (
            O => \N__23126\,
            I => \N__23122\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__23125\,
            I => \N__23119\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__23122\,
            I => \N__23116\
        );

    \I__2272\ : InMux
    port map (
            O => \N__23119\,
            I => \N__23113\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__23116\,
            I => \pwm_generator_inst.un18_threshold1_18\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__23113\,
            I => \pwm_generator_inst.un18_threshold1_18\
        );

    \I__2269\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23105\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__23105\,
            I => \N__23102\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__23102\,
            I => \pwm_generator_inst.un22_threshold_1_cry_0_THRU_CO\
        );

    \I__2266\ : InMux
    port map (
            O => \N__23099\,
            I => \pwm_generator_inst.un22_threshold_1_cry_0\
        );

    \I__2265\ : InMux
    port map (
            O => \N__23096\,
            I => \pwm_generator_inst.un22_threshold_1_cry_1\
        );

    \I__2264\ : InMux
    port map (
            O => \N__23093\,
            I => \pwm_generator_inst.un22_threshold_1_cry_2\
        );

    \I__2263\ : InMux
    port map (
            O => \N__23090\,
            I => \pwm_generator_inst.un22_threshold_1_cry_3\
        );

    \I__2262\ : InMux
    port map (
            O => \N__23087\,
            I => \pwm_generator_inst.un22_threshold_1_cry_4\
        );

    \I__2261\ : InMux
    port map (
            O => \N__23084\,
            I => \pwm_generator_inst.un22_threshold_1_cry_5\
        );

    \I__2260\ : InMux
    port map (
            O => \N__23081\,
            I => \pwm_generator_inst.un22_threshold_1_cry_6\
        );

    \I__2259\ : InMux
    port map (
            O => \N__23078\,
            I => \pwm_generator_inst.un3_threshold_cry_16\
        );

    \I__2258\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23072\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__23072\,
            I => \N__23069\
        );

    \I__2256\ : Span4Mux_s1_h
    port map (
            O => \N__23069\,
            I => \N__23066\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__23066\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFDZ0\
        );

    \I__2254\ : InMux
    port map (
            O => \N__23063\,
            I => \pwm_generator_inst.un3_threshold_cry_17\
        );

    \I__2253\ : InMux
    port map (
            O => \N__23060\,
            I => \pwm_generator_inst.un3_threshold_cry_18\
        );

    \I__2252\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23054\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__23054\,
            I => \N__23051\
        );

    \I__2250\ : Span4Mux_v
    port map (
            O => \N__23051\,
            I => \N__23048\
        );

    \I__2249\ : Odrv4
    port map (
            O => \N__23048\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__2248\ : InMux
    port map (
            O => \N__23045\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__23042\,
            I => \N__23039\
        );

    \I__2246\ : InMux
    port map (
            O => \N__23039\,
            I => \N__23036\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__23036\,
            I => \N__23033\
        );

    \I__2244\ : Span4Mux_v
    port map (
            O => \N__23033\,
            I => \N__23030\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__23030\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNOZ0\
        );

    \I__2242\ : InMux
    port map (
            O => \N__23027\,
            I => \N__23024\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__23024\,
            I => \N_112_i_i\
        );

    \I__2240\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23018\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__23018\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__23015\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__2237\ : InMux
    port map (
            O => \N__23012\,
            I => \N__23009\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__23009\,
            I => \N__23006\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__23006\,
            I => \N__23002\
        );

    \I__2234\ : InMux
    port map (
            O => \N__23005\,
            I => \N__22999\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__23002\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__22999\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0\
        );

    \I__2231\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22991\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__22991\,
            I => \N__22988\
        );

    \I__2229\ : Span4Mux_v
    port map (
            O => \N__22988\,
            I => \N__22985\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__22985\,
            I => \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDIZ0Z8\
        );

    \I__2227\ : InMux
    port map (
            O => \N__22982\,
            I => \pwm_generator_inst.un3_threshold_cry_8\
        );

    \I__2226\ : InMux
    port map (
            O => \N__22979\,
            I => \N__22976\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__22976\,
            I => \N__22973\
        );

    \I__2224\ : Span4Mux_v
    port map (
            O => \N__22973\,
            I => \N__22970\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__22970\,
            I => \pwm_generator_inst.un3_threshold_cry_9_c_RNISHKZ0Z8\
        );

    \I__2222\ : InMux
    port map (
            O => \N__22967\,
            I => \pwm_generator_inst.un3_threshold_cry_9\
        );

    \I__2221\ : InMux
    port map (
            O => \N__22964\,
            I => \N__22961\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__22961\,
            I => \N__22958\
        );

    \I__2219\ : Span4Mux_v
    port map (
            O => \N__22958\,
            I => \N__22955\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__22955\,
            I => \pwm_generator_inst.un3_threshold_cry_10_c_RNI59GZ0Z7\
        );

    \I__2217\ : InMux
    port map (
            O => \N__22952\,
            I => \pwm_generator_inst.un3_threshold_cry_10\
        );

    \I__2216\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22946\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__22946\,
            I => \N__22943\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__22943\,
            I => \N__22940\
        );

    \I__2213\ : Odrv4
    port map (
            O => \N__22940\,
            I => \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DIZ0Z7\
        );

    \I__2212\ : InMux
    port map (
            O => \N__22937\,
            I => \pwm_generator_inst.un3_threshold_cry_11\
        );

    \I__2211\ : InMux
    port map (
            O => \N__22934\,
            I => \N__22931\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__22931\,
            I => \N__22928\
        );

    \I__2209\ : Span4Mux_v
    port map (
            O => \N__22928\,
            I => \N__22925\
        );

    \I__2208\ : Odrv4
    port map (
            O => \N__22925\,
            I => \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HKZ0Z7\
        );

    \I__2207\ : InMux
    port map (
            O => \N__22922\,
            I => \pwm_generator_inst.un3_threshold_cry_12\
        );

    \I__2206\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22916\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__22916\,
            I => \N__22913\
        );

    \I__2204\ : Span4Mux_v
    port map (
            O => \N__22913\,
            I => \N__22910\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__22910\,
            I => \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLMZ0Z7\
        );

    \I__2202\ : InMux
    port map (
            O => \N__22907\,
            I => \pwm_generator_inst.un3_threshold_cry_13\
        );

    \I__2201\ : InMux
    port map (
            O => \N__22904\,
            I => \N__22901\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__22901\,
            I => \N__22898\
        );

    \I__2199\ : Span4Mux_v
    port map (
            O => \N__22898\,
            I => \N__22895\
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__22895\,
            I => \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPOZ0Z7\
        );

    \I__2197\ : InMux
    port map (
            O => \N__22892\,
            I => \pwm_generator_inst.un3_threshold_cry_14\
        );

    \I__2196\ : InMux
    port map (
            O => \N__22889\,
            I => \N__22886\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__22886\,
            I => \N__22883\
        );

    \I__2194\ : Span4Mux_v
    port map (
            O => \N__22883\,
            I => \N__22880\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__22880\,
            I => \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQZ0Z7\
        );

    \I__2192\ : InMux
    port map (
            O => \N__22877\,
            I => \bfn_1_22_0_\
        );

    \I__2191\ : InMux
    port map (
            O => \N__22874\,
            I => \N__22871\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__22871\,
            I => \N__22868\
        );

    \I__2189\ : Span4Mux_v
    port map (
            O => \N__22868\,
            I => \N__22865\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__22865\,
            I => \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1TZ0Z7\
        );

    \I__2187\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22859\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__22859\,
            I => \N__22856\
        );

    \I__2185\ : Span12Mux_v
    port map (
            O => \N__22856\,
            I => \N__22853\
        );

    \I__2184\ : Span12Mux_h
    port map (
            O => \N__22853\,
            I => \N__22850\
        );

    \I__2183\ : Span12Mux_h
    port map (
            O => \N__22850\,
            I => \N__22847\
        );

    \I__2182\ : Odrv12
    port map (
            O => \N__22847\,
            I => \pwm_generator_inst.O_0_8\
        );

    \I__2181\ : InMux
    port map (
            O => \N__22844\,
            I => \N__22841\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__22841\,
            I => \N__22838\
        );

    \I__2179\ : Span4Mux_v
    port map (
            O => \N__22838\,
            I => \N__22835\
        );

    \I__2178\ : Sp12to4
    port map (
            O => \N__22835\,
            I => \N__22832\
        );

    \I__2177\ : Odrv12
    port map (
            O => \N__22832\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CCZ0\
        );

    \I__2176\ : InMux
    port map (
            O => \N__22829\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__22826\,
            I => \N__22823\
        );

    \I__2174\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22820\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__22820\,
            I => \N__22817\
        );

    \I__2172\ : Span12Mux_v
    port map (
            O => \N__22817\,
            I => \N__22814\
        );

    \I__2171\ : Span12Mux_h
    port map (
            O => \N__22814\,
            I => \N__22811\
        );

    \I__2170\ : Span12Mux_h
    port map (
            O => \N__22811\,
            I => \N__22808\
        );

    \I__2169\ : Odrv12
    port map (
            O => \N__22808\,
            I => \pwm_generator_inst.O_0_9\
        );

    \I__2168\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22802\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__22802\,
            I => \N__22799\
        );

    \I__2166\ : Span4Mux_v
    port map (
            O => \N__22799\,
            I => \N__22796\
        );

    \I__2165\ : Sp12to4
    port map (
            O => \N__22796\,
            I => \N__22793\
        );

    \I__2164\ : Odrv12
    port map (
            O => \N__22793\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DCZ0\
        );

    \I__2163\ : InMux
    port map (
            O => \N__22790\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__2162\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22784\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__22784\,
            I => \N__22781\
        );

    \I__2160\ : Span12Mux_v
    port map (
            O => \N__22781\,
            I => \N__22778\
        );

    \I__2159\ : Span12Mux_h
    port map (
            O => \N__22778\,
            I => \N__22775\
        );

    \I__2158\ : Span12Mux_h
    port map (
            O => \N__22775\,
            I => \N__22772\
        );

    \I__2157\ : Odrv12
    port map (
            O => \N__22772\,
            I => \pwm_generator_inst.O_0_10\
        );

    \I__2156\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22766\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__22766\,
            I => \N__22763\
        );

    \I__2154\ : Span12Mux_s1_h
    port map (
            O => \N__22763\,
            I => \N__22760\
        );

    \I__2153\ : Span12Mux_v
    port map (
            O => \N__22760\,
            I => \N__22757\
        );

    \I__2152\ : Odrv12
    port map (
            O => \N__22757\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI77ECZ0\
        );

    \I__2151\ : InMux
    port map (
            O => \N__22754\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__2150\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22748\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__22748\,
            I => \N__22745\
        );

    \I__2148\ : Span12Mux_v
    port map (
            O => \N__22745\,
            I => \N__22742\
        );

    \I__2147\ : Span12Mux_h
    port map (
            O => \N__22742\,
            I => \N__22739\
        );

    \I__2146\ : Span12Mux_h
    port map (
            O => \N__22739\,
            I => \N__22736\
        );

    \I__2145\ : Odrv12
    port map (
            O => \N__22736\,
            I => \pwm_generator_inst.O_0_11\
        );

    \I__2144\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22730\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__22730\,
            I => \N__22727\
        );

    \I__2142\ : Span4Mux_v
    port map (
            O => \N__22727\,
            I => \N__22724\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__22724\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FCZ0\
        );

    \I__2140\ : InMux
    port map (
            O => \N__22721\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__2139\ : InMux
    port map (
            O => \N__22718\,
            I => \N__22715\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__22715\,
            I => \N__22712\
        );

    \I__2137\ : Span12Mux_h
    port map (
            O => \N__22712\,
            I => \N__22709\
        );

    \I__2136\ : Span12Mux_h
    port map (
            O => \N__22709\,
            I => \N__22706\
        );

    \I__2135\ : Odrv12
    port map (
            O => \N__22706\,
            I => \pwm_generator_inst.O_0_12\
        );

    \I__2134\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22700\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__22700\,
            I => \N__22697\
        );

    \I__2132\ : Span4Mux_v
    port map (
            O => \N__22697\,
            I => \N__22694\
        );

    \I__2131\ : Odrv4
    port map (
            O => \N__22694\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGCZ0\
        );

    \I__2130\ : InMux
    port map (
            O => \N__22691\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__2129\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22685\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__22685\,
            I => \N__22682\
        );

    \I__2127\ : Span4Mux_v
    port map (
            O => \N__22682\,
            I => \N__22679\
        );

    \I__2126\ : Sp12to4
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__2125\ : Span12Mux_h
    port map (
            O => \N__22676\,
            I => \N__22673\
        );

    \I__2124\ : Span12Mux_h
    port map (
            O => \N__22673\,
            I => \N__22670\
        );

    \I__2123\ : Odrv12
    port map (
            O => \N__22670\,
            I => \pwm_generator_inst.O_0_13\
        );

    \I__2122\ : InMux
    port map (
            O => \N__22667\,
            I => \N__22664\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__22664\,
            I => \N__22661\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__22661\,
            I => \N__22658\
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__22658\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHCZ0\
        );

    \I__2118\ : InMux
    port map (
            O => \N__22655\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__2117\ : InMux
    port map (
            O => \N__22652\,
            I => \N__22649\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__22649\,
            I => \N__22646\
        );

    \I__2115\ : Span4Mux_v
    port map (
            O => \N__22646\,
            I => \N__22643\
        );

    \I__2114\ : Sp12to4
    port map (
            O => \N__22643\,
            I => \N__22640\
        );

    \I__2113\ : Span12Mux_h
    port map (
            O => \N__22640\,
            I => \N__22637\
        );

    \I__2112\ : Odrv12
    port map (
            O => \N__22637\,
            I => \pwm_generator_inst.O_0_14\
        );

    \I__2111\ : InMux
    port map (
            O => \N__22634\,
            I => \N__22631\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__22631\,
            I => \N__22628\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__22628\,
            I => \N__22625\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__22625\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFICZ0\
        );

    \I__2107\ : InMux
    port map (
            O => \N__22622\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__2106\ : InMux
    port map (
            O => \N__22619\,
            I => \N__22616\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__22616\,
            I => \N__22613\
        );

    \I__2104\ : Span4Mux_v
    port map (
            O => \N__22613\,
            I => \N__22610\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__22610\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FOZ0\
        );

    \I__2102\ : InMux
    port map (
            O => \N__22607\,
            I => \bfn_1_21_0_\
        );

    \I__2101\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22601\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22598\
        );

    \I__2099\ : Span4Mux_v
    port map (
            O => \N__22598\,
            I => \N__22595\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__22595\,
            I => \N__22592\
        );

    \I__2097\ : Odrv4
    port map (
            O => \N__22592\,
            I => \pwm_generator_inst.un5_threshold_1_25\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__22589\,
            I => \N__22586\
        );

    \I__2095\ : InMux
    port map (
            O => \N__22586\,
            I => \N__22583\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__22583\,
            I => \N__22580\
        );

    \I__2093\ : Span4Mux_v
    port map (
            O => \N__22580\,
            I => \N__22577\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__22577\,
            I => \pwm_generator_inst.un5_threshold_2_10\
        );

    \I__2091\ : InMux
    port map (
            O => \N__22574\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_9\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__22571\,
            I => \N__22568\
        );

    \I__2089\ : InMux
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__22565\,
            I => \N__22562\
        );

    \I__2087\ : Span4Mux_v
    port map (
            O => \N__22562\,
            I => \N__22559\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__22559\,
            I => \pwm_generator_inst.un5_threshold_2_11\
        );

    \I__2085\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22553\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__22550\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPFZ0\
        );

    \I__2082\ : InMux
    port map (
            O => \N__22547\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_10\
        );

    \I__2081\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22541\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__22541\,
            I => \N__22538\
        );

    \I__2079\ : Span4Mux_v
    port map (
            O => \N__22538\,
            I => \N__22535\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__22535\,
            I => \pwm_generator_inst.un5_threshold_2_12\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__22532\,
            I => \N__22529\
        );

    \I__2076\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22526\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__22526\,
            I => \N__22523\
        );

    \I__2074\ : Span4Mux_v
    port map (
            O => \N__22523\,
            I => \N__22520\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__22520\,
            I => \pwm_generator_inst.un5_threshold_2_13\
        );

    \I__2072\ : InMux
    port map (
            O => \N__22517\,
            I => \N__22514\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__22514\,
            I => \N__22511\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__22511\,
            I => \N__22508\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__22508\,
            I => \pwm_generator_inst.un5_threshold_2_14\
        );

    \I__2068\ : InMux
    port map (
            O => \N__22505\,
            I => \bfn_1_19_0_\
        );

    \I__2067\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22499\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__2065\ : Span4Mux_v
    port map (
            O => \N__22496\,
            I => \N__22493\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__22493\,
            I => \pwm_generator_inst.un5_threshold_2_2\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__22490\,
            I => \N__22487\
        );

    \I__2062\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22484\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__22484\,
            I => \N__22481\
        );

    \I__2060\ : Span4Mux_v
    port map (
            O => \N__22481\,
            I => \N__22478\
        );

    \I__2059\ : Span4Mux_v
    port map (
            O => \N__22478\,
            I => \N__22475\
        );

    \I__2058\ : Odrv4
    port map (
            O => \N__22475\,
            I => \pwm_generator_inst.un5_threshold_1_17\
        );

    \I__2057\ : InMux
    port map (
            O => \N__22472\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_1\
        );

    \I__2056\ : InMux
    port map (
            O => \N__22469\,
            I => \N__22466\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__22466\,
            I => \N__22463\
        );

    \I__2054\ : Span4Mux_v
    port map (
            O => \N__22463\,
            I => \N__22460\
        );

    \I__2053\ : Odrv4
    port map (
            O => \N__22460\,
            I => \pwm_generator_inst.un5_threshold_2_3\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__22457\,
            I => \N__22454\
        );

    \I__2051\ : InMux
    port map (
            O => \N__22454\,
            I => \N__22451\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__22451\,
            I => \N__22448\
        );

    \I__2049\ : Span4Mux_v
    port map (
            O => \N__22448\,
            I => \N__22445\
        );

    \I__2048\ : Span4Mux_s1_h
    port map (
            O => \N__22445\,
            I => \N__22442\
        );

    \I__2047\ : Span4Mux_v
    port map (
            O => \N__22442\,
            I => \N__22439\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__22439\,
            I => \pwm_generator_inst.un5_threshold_1_18\
        );

    \I__2045\ : InMux
    port map (
            O => \N__22436\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_2\
        );

    \I__2044\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22430\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__22430\,
            I => \N__22427\
        );

    \I__2042\ : Span4Mux_v
    port map (
            O => \N__22427\,
            I => \N__22424\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__22424\,
            I => \pwm_generator_inst.un5_threshold_2_4\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__22421\,
            I => \N__22418\
        );

    \I__2039\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22415\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__22415\,
            I => \N__22412\
        );

    \I__2037\ : Span4Mux_v
    port map (
            O => \N__22412\,
            I => \N__22409\
        );

    \I__2036\ : Span4Mux_v
    port map (
            O => \N__22409\,
            I => \N__22406\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__22406\,
            I => \pwm_generator_inst.un5_threshold_1_19\
        );

    \I__2034\ : InMux
    port map (
            O => \N__22403\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_3\
        );

    \I__2033\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22397\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__22397\,
            I => \N__22394\
        );

    \I__2031\ : Span4Mux_v
    port map (
            O => \N__22394\,
            I => \N__22391\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__22391\,
            I => \pwm_generator_inst.un5_threshold_2_5\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__22388\,
            I => \N__22385\
        );

    \I__2028\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22382\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__22382\,
            I => \N__22379\
        );

    \I__2026\ : Span4Mux_v
    port map (
            O => \N__22379\,
            I => \N__22376\
        );

    \I__2025\ : Span4Mux_v
    port map (
            O => \N__22376\,
            I => \N__22373\
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__22373\,
            I => \pwm_generator_inst.un5_threshold_1_20\
        );

    \I__2023\ : InMux
    port map (
            O => \N__22370\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_4\
        );

    \I__2022\ : InMux
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__22364\,
            I => \N__22361\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__22361\,
            I => \N__22358\
        );

    \I__2019\ : Span4Mux_v
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__22355\,
            I => \pwm_generator_inst.un5_threshold_1_21\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__2016\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__22340\,
            I => \pwm_generator_inst.un5_threshold_2_6\
        );

    \I__2012\ : InMux
    port map (
            O => \N__22337\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_5\
        );

    \I__2011\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__22331\,
            I => \N__22328\
        );

    \I__2009\ : Span4Mux_v
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__2008\ : Span4Mux_v
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__22322\,
            I => \pwm_generator_inst.un5_threshold_1_22\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__22319\,
            I => \N__22316\
        );

    \I__2005\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__22307\,
            I => \pwm_generator_inst.un5_threshold_2_7\
        );

    \I__2001\ : InMux
    port map (
            O => \N__22304\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_6\
        );

    \I__2000\ : InMux
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__1998\ : Span4Mux_v
    port map (
            O => \N__22295\,
            I => \N__22292\
        );

    \I__1997\ : Span4Mux_v
    port map (
            O => \N__22292\,
            I => \N__22289\
        );

    \I__1996\ : Odrv4
    port map (
            O => \N__22289\,
            I => \pwm_generator_inst.un5_threshold_1_23\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__22286\,
            I => \N__22283\
        );

    \I__1994\ : InMux
    port map (
            O => \N__22283\,
            I => \N__22280\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__22280\,
            I => \N__22277\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__22274\,
            I => \pwm_generator_inst.un5_threshold_2_8\
        );

    \I__1990\ : InMux
    port map (
            O => \N__22271\,
            I => \bfn_1_18_0_\
        );

    \I__1989\ : InMux
    port map (
            O => \N__22268\,
            I => \N__22265\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__22265\,
            I => \N__22262\
        );

    \I__1987\ : Span4Mux_v
    port map (
            O => \N__22262\,
            I => \N__22259\
        );

    \I__1986\ : Span4Mux_v
    port map (
            O => \N__22259\,
            I => \N__22256\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__22256\,
            I => \pwm_generator_inst.un5_threshold_1_24\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__22253\,
            I => \N__22250\
        );

    \I__1983\ : InMux
    port map (
            O => \N__22250\,
            I => \N__22247\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__22247\,
            I => \N__22244\
        );

    \I__1981\ : Span4Mux_v
    port map (
            O => \N__22244\,
            I => \N__22241\
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__22241\,
            I => \pwm_generator_inst.un5_threshold_2_9\
        );

    \I__1979\ : InMux
    port map (
            O => \N__22238\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_8\
        );

    \I__1978\ : InMux
    port map (
            O => \N__22235\,
            I => \pwm_generator_inst.un18_threshold_1_cry_24\
        );

    \I__1977\ : InMux
    port map (
            O => \N__22232\,
            I => \pwm_generator_inst.un18_threshold_1_cry_25\
        );

    \I__1976\ : InMux
    port map (
            O => \N__22229\,
            I => \N__22226\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__22226\,
            I => \pwm_generator_inst.un18_threshold_1_axb_20\
        );

    \I__1974\ : InMux
    port map (
            O => \N__22223\,
            I => \N__22220\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__22220\,
            I => \pwm_generator_inst.un18_threshold_1_axb_17\
        );

    \I__1972\ : InMux
    port map (
            O => \N__22217\,
            I => \N__22214\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__22214\,
            I => \pwm_generator_inst.un18_threshold_1_axb_18\
        );

    \I__1970\ : InMux
    port map (
            O => \N__22211\,
            I => \N__22208\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__22208\,
            I => \pwm_generator_inst.un18_threshold_1_axb_22\
        );

    \I__1968\ : InMux
    port map (
            O => \N__22205\,
            I => \N__22202\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__22202\,
            I => \pwm_generator_inst.un18_threshold_1_axb_21\
        );

    \I__1966\ : InMux
    port map (
            O => \N__22199\,
            I => \N__22196\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__1964\ : Span4Mux_v
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__22190\,
            I => \pwm_generator_inst.un5_threshold_2_0\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__1961\ : InMux
    port map (
            O => \N__22184\,
            I => \N__22181\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__1959\ : Span12Mux_v
    port map (
            O => \N__22178\,
            I => \N__22175\
        );

    \I__1958\ : Odrv12
    port map (
            O => \N__22175\,
            I => \pwm_generator_inst.un5_threshold_1_15\
        );

    \I__1957\ : InMux
    port map (
            O => \N__22172\,
            I => \N__22169\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__1955\ : Odrv4
    port map (
            O => \N__22166\,
            I => \pwm_generator_inst.un18_threshold_1_axb_15\
        );

    \I__1954\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22160\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__22160\,
            I => \N__22157\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__22157\,
            I => \N__22154\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__22154\,
            I => \pwm_generator_inst.un5_threshold_2_1\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__22151\,
            I => \N__22148\
        );

    \I__1949\ : InMux
    port map (
            O => \N__22148\,
            I => \N__22145\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__1946\ : Span4Mux_v
    port map (
            O => \N__22139\,
            I => \N__22136\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__22136\,
            I => \pwm_generator_inst.un5_threshold_1_16\
        );

    \I__1944\ : InMux
    port map (
            O => \N__22133\,
            I => \N__22130\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__22130\,
            I => \N__22127\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__22127\,
            I => \pwm_generator_inst.un18_threshold_1_axb_16\
        );

    \I__1941\ : InMux
    port map (
            O => \N__22124\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_0\
        );

    \I__1940\ : InMux
    port map (
            O => \N__22121\,
            I => \pwm_generator_inst.un18_threshold_1_cry_16\
        );

    \I__1939\ : InMux
    port map (
            O => \N__22118\,
            I => \pwm_generator_inst.un18_threshold_1_cry_17\
        );

    \I__1938\ : InMux
    port map (
            O => \N__22115\,
            I => \pwm_generator_inst.un18_threshold_1_cry_18\
        );

    \I__1937\ : InMux
    port map (
            O => \N__22112\,
            I => \pwm_generator_inst.un18_threshold_1_cry_19\
        );

    \I__1936\ : InMux
    port map (
            O => \N__22109\,
            I => \pwm_generator_inst.un18_threshold_1_cry_20\
        );

    \I__1935\ : InMux
    port map (
            O => \N__22106\,
            I => \pwm_generator_inst.un18_threshold_1_cry_21\
        );

    \I__1934\ : InMux
    port map (
            O => \N__22103\,
            I => \pwm_generator_inst.un18_threshold_1_cry_22\
        );

    \I__1933\ : InMux
    port map (
            O => \N__22100\,
            I => \bfn_1_16_0_\
        );

    \I__1932\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22094\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__22094\,
            I => \N__22091\
        );

    \I__1930\ : Span12Mux_h
    port map (
            O => \N__22091\,
            I => \N__22088\
        );

    \I__1929\ : Odrv12
    port map (
            O => \N__22088\,
            I => \pwm_generator_inst.O_8\
        );

    \I__1928\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22082\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__22082\,
            I => \pwm_generator_inst.un18_threshold_1_axb_8\
        );

    \I__1926\ : InMux
    port map (
            O => \N__22079\,
            I => \N__22076\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__22076\,
            I => \N__22073\
        );

    \I__1924\ : Span4Mux_v
    port map (
            O => \N__22073\,
            I => \N__22070\
        );

    \I__1923\ : Span4Mux_v
    port map (
            O => \N__22070\,
            I => \N__22067\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__22067\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1921\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22061\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__22061\,
            I => \pwm_generator_inst.un18_threshold_1_axb_9\
        );

    \I__1919\ : InMux
    port map (
            O => \N__22058\,
            I => \N__22055\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__22055\,
            I => \N__22052\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__22052\,
            I => \N__22049\
        );

    \I__1916\ : Span4Mux_v
    port map (
            O => \N__22049\,
            I => \N__22046\
        );

    \I__1915\ : Odrv4
    port map (
            O => \N__22046\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1914\ : InMux
    port map (
            O => \N__22043\,
            I => \N__22040\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__22040\,
            I => \pwm_generator_inst.un18_threshold_1_axb_10\
        );

    \I__1912\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22034\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__22034\,
            I => \N__22031\
        );

    \I__1910\ : Span4Mux_v
    port map (
            O => \N__22031\,
            I => \N__22028\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__22028\,
            I => \N__22025\
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__22025\,
            I => \pwm_generator_inst.O_11\
        );

    \I__1907\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22019\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__22019\,
            I => \pwm_generator_inst.un18_threshold_1_axb_11\
        );

    \I__1905\ : InMux
    port map (
            O => \N__22016\,
            I => \N__22013\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__22013\,
            I => \N__22010\
        );

    \I__1903\ : Span4Mux_v
    port map (
            O => \N__22010\,
            I => \N__22007\
        );

    \I__1902\ : Span4Mux_v
    port map (
            O => \N__22007\,
            I => \N__22004\
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__22004\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1900\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__21998\,
            I => \pwm_generator_inst.un18_threshold_1_axb_12\
        );

    \I__1898\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21992\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__21992\,
            I => \N__21989\
        );

    \I__1896\ : Span4Mux_v
    port map (
            O => \N__21989\,
            I => \N__21986\
        );

    \I__1895\ : Span4Mux_v
    port map (
            O => \N__21986\,
            I => \N__21983\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__21983\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1893\ : InMux
    port map (
            O => \N__21980\,
            I => \N__21977\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__21977\,
            I => \pwm_generator_inst.un18_threshold_1_axb_13\
        );

    \I__1891\ : InMux
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__21971\,
            I => \N__21968\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__21968\,
            I => \N__21965\
        );

    \I__1888\ : Span4Mux_v
    port map (
            O => \N__21965\,
            I => \N__21962\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__21962\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1886\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21956\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__21956\,
            I => \pwm_generator_inst.un18_threshold_1_axb_14\
        );

    \I__1884\ : InMux
    port map (
            O => \N__21953\,
            I => \N__21950\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__1882\ : Span4Mux_v
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__1881\ : Span4Mux_v
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__21941\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1879\ : InMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__21935\,
            I => \pwm_generator_inst.un18_threshold_1_axb_1\
        );

    \I__1877\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__21926\,
            I => \N__21923\
        );

    \I__1874\ : Span4Mux_v
    port map (
            O => \N__21923\,
            I => \N__21920\
        );

    \I__1873\ : Odrv4
    port map (
            O => \N__21920\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1872\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21914\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__21914\,
            I => \pwm_generator_inst.un18_threshold_1_axb_2\
        );

    \I__1870\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21908\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__21908\,
            I => \N__21905\
        );

    \I__1868\ : Span4Mux_v
    port map (
            O => \N__21905\,
            I => \N__21902\
        );

    \I__1867\ : Span4Mux_v
    port map (
            O => \N__21902\,
            I => \N__21899\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__21899\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1865\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21893\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__21893\,
            I => \pwm_generator_inst.un18_threshold_1_axb_3\
        );

    \I__1863\ : InMux
    port map (
            O => \N__21890\,
            I => \N__21887\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__21887\,
            I => \N__21884\
        );

    \I__1861\ : Span4Mux_v
    port map (
            O => \N__21884\,
            I => \N__21881\
        );

    \I__1860\ : Span4Mux_v
    port map (
            O => \N__21881\,
            I => \N__21878\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__21878\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1858\ : InMux
    port map (
            O => \N__21875\,
            I => \N__21872\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__21872\,
            I => \pwm_generator_inst.un18_threshold_1_axb_4\
        );

    \I__1856\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21866\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__21866\,
            I => \N__21863\
        );

    \I__1854\ : Span4Mux_v
    port map (
            O => \N__21863\,
            I => \N__21860\
        );

    \I__1853\ : Span4Mux_v
    port map (
            O => \N__21860\,
            I => \N__21857\
        );

    \I__1852\ : Odrv4
    port map (
            O => \N__21857\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1851\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21851\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__21851\,
            I => \pwm_generator_inst.un18_threshold_1_axb_5\
        );

    \I__1849\ : InMux
    port map (
            O => \N__21848\,
            I => \N__21845\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__21845\,
            I => \N__21842\
        );

    \I__1847\ : Span4Mux_v
    port map (
            O => \N__21842\,
            I => \N__21839\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__21839\,
            I => \N__21836\
        );

    \I__1845\ : Odrv4
    port map (
            O => \N__21836\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1844\ : InMux
    port map (
            O => \N__21833\,
            I => \N__21830\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__21830\,
            I => \pwm_generator_inst.un18_threshold_1_axb_6\
        );

    \I__1842\ : InMux
    port map (
            O => \N__21827\,
            I => \N__21824\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__21824\,
            I => \N__21821\
        );

    \I__1840\ : Span12Mux_v
    port map (
            O => \N__21821\,
            I => \N__21818\
        );

    \I__1839\ : Odrv12
    port map (
            O => \N__21818\,
            I => \pwm_generator_inst.O_7\
        );

    \I__1838\ : InMux
    port map (
            O => \N__21815\,
            I => \N__21812\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__21812\,
            I => \pwm_generator_inst.un18_threshold_1_axb_7\
        );

    \I__1836\ : InMux
    port map (
            O => \N__21809\,
            I => \N__21806\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__21806\,
            I => \N__21803\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__21803\,
            I => \N__21800\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__21797\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1831\ : InMux
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__21791\,
            I => \pwm_generator_inst.un18_threshold_1_axb_0\
        );

    \I__1829\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__1827\ : Sp12to4
    port map (
            O => \N__21782\,
            I => \N__21779\
        );

    \I__1826\ : Span12Mux_s11_v
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__1825\ : Span12Mux_h
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__1824\ : Span12Mux_h
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__1823\ : Odrv12
    port map (
            O => \N__21770\,
            I => \pwm_generator_inst.O_0_1\
        );

    \I__1822\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__1820\ : Sp12to4
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__1819\ : Span12Mux_s10_v
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__1818\ : Span12Mux_h
    port map (
            O => \N__21755\,
            I => \N__21752\
        );

    \I__1817\ : Span12Mux_h
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__1816\ : Odrv12
    port map (
            O => \N__21749\,
            I => \pwm_generator_inst.O_0_0\
        );

    \I__1815\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21743\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__21743\,
            I => \N__21740\
        );

    \I__1813\ : Span4Mux_v
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__1812\ : Sp12to4
    port map (
            O => \N__21737\,
            I => \N__21734\
        );

    \I__1811\ : Span12Mux_h
    port map (
            O => \N__21734\,
            I => \N__21731\
        );

    \I__1810\ : Span12Mux_h
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__1809\ : Span12Mux_v
    port map (
            O => \N__21728\,
            I => \N__21725\
        );

    \I__1808\ : Odrv12
    port map (
            O => \N__21725\,
            I => \pwm_generator_inst.O_0_5\
        );

    \I__1807\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21719\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__21719\,
            I => \N__21716\
        );

    \I__1805\ : Sp12to4
    port map (
            O => \N__21716\,
            I => \N__21713\
        );

    \I__1804\ : Span12Mux_s5_v
    port map (
            O => \N__21713\,
            I => \N__21710\
        );

    \I__1803\ : Span12Mux_h
    port map (
            O => \N__21710\,
            I => \N__21707\
        );

    \I__1802\ : Span12Mux_h
    port map (
            O => \N__21707\,
            I => \N__21704\
        );

    \I__1801\ : Odrv12
    port map (
            O => \N__21704\,
            I => \pwm_generator_inst.O_0_3\
        );

    \I__1800\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21698\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__21698\,
            I => \N__21695\
        );

    \I__1798\ : Span12Mux_s1_h
    port map (
            O => \N__21695\,
            I => \N__21692\
        );

    \I__1797\ : Span12Mux_h
    port map (
            O => \N__21692\,
            I => \N__21689\
        );

    \I__1796\ : Span12Mux_h
    port map (
            O => \N__21689\,
            I => \N__21686\
        );

    \I__1795\ : Odrv12
    port map (
            O => \N__21686\,
            I => \pwm_generator_inst.O_0_4\
        );

    \I__1794\ : InMux
    port map (
            O => \N__21683\,
            I => \N__21680\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__1792\ : Sp12to4
    port map (
            O => \N__21677\,
            I => \N__21674\
        );

    \I__1791\ : Span12Mux_v
    port map (
            O => \N__21674\,
            I => \N__21671\
        );

    \I__1790\ : Span12Mux_h
    port map (
            O => \N__21671\,
            I => \N__21668\
        );

    \I__1789\ : Span12Mux_h
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__1788\ : Odrv12
    port map (
            O => \N__21665\,
            I => \pwm_generator_inst.O_0_2\
        );

    \I__1787\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21659\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__21659\,
            I => \N__21656\
        );

    \I__1785\ : Span4Mux_v
    port map (
            O => \N__21656\,
            I => \N__21653\
        );

    \I__1784\ : Sp12to4
    port map (
            O => \N__21653\,
            I => \N__21650\
        );

    \I__1783\ : Span12Mux_h
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__1782\ : Span12Mux_h
    port map (
            O => \N__21647\,
            I => \N__21644\
        );

    \I__1781\ : Odrv12
    port map (
            O => \N__21644\,
            I => \pwm_generator_inst.O_0_6\
        );

    \I__1780\ : IoInMux
    port map (
            O => \N__21641\,
            I => \N__21638\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__21638\,
            I => \N__21635\
        );

    \I__1778\ : IoSpan4Mux
    port map (
            O => \N__21635\,
            I => \N__21632\
        );

    \I__1777\ : IoSpan4Mux
    port map (
            O => \N__21632\,
            I => \N__21629\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__21629\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \I__1775\ : IoInMux
    port map (
            O => \N__21626\,
            I => \N__21623\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__21623\,
            I => \N__21620\
        );

    \I__1773\ : Span4Mux_s3_v
    port map (
            O => \N__21620\,
            I => \N__21617\
        );

    \I__1772\ : Span4Mux_h
    port map (
            O => \N__21617\,
            I => \N__21614\
        );

    \I__1771\ : Sp12to4
    port map (
            O => \N__21614\,
            I => \N__21611\
        );

    \I__1770\ : Span12Mux_v
    port map (
            O => \N__21611\,
            I => \N__21608\
        );

    \I__1769\ : Span12Mux_v
    port map (
            O => \N__21608\,
            I => \N__21605\
        );

    \I__1768\ : Odrv12
    port map (
            O => \N__21605\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_1_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_20_0_\
        );

    \IN_MUX_bfv_1_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_1_21_0_\
        );

    \IN_MUX_bfv_1_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_1_22_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un22_threshold_1_cry_7\,
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_16_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_13_0_\
        );

    \IN_MUX_bfv_16_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_16_14_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_18_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_23_0_\
        );

    \IN_MUX_bfv_18_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryinitout => \bfn_18_24_0_\
        );

    \IN_MUX_bfv_18_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryinitout => \bfn_18_25_0_\
        );

    \IN_MUX_bfv_18_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryinitout => \bfn_18_26_0_\
        );

    \IN_MUX_bfv_13_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_21_0_\
        );

    \IN_MUX_bfv_13_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_13_22_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un5_threshold_add_1_cry_7\,
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un5_threshold_add_1_cry_15\,
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un18_threshold_1_cry_7\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un18_threshold_1_cry_15\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un18_threshold_1_cry_23\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_3_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_15_0_\
        );

    \IN_MUX_bfv_3_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_3_16_0_\
        );

    \IN_MUX_bfv_3_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_12_0_\
        );

    \IN_MUX_bfv_3_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_3_13_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_7\,
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_15\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_30\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.counter_cry_7\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.counter_cry_15\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.counter_cry_23\,
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_11_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_4_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_7\,
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_15\,
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_30\,
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_10_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_2_0_\
        );

    \IN_MUX_bfv_10_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.counter_cry_7\,
            carryinitout => \bfn_10_3_0_\
        );

    \IN_MUX_bfv_10_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.counter_cry_15\,
            carryinitout => \bfn_10_4_0_\
        );

    \IN_MUX_bfv_10_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.counter_cry_23\,
            carryinitout => \bfn_10_5_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_7\,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_15\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_30\,
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16\,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24\,
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7\,
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23\,
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.counter_cry_7\,
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_8_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.counter_cry_15\,
            carryinitout => \bfn_8_22_0_\
        );

    \IN_MUX_bfv_8_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.counter_cry_23\,
            carryinitout => \bfn_8_23_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_7\,
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_15\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_30\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8\,
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16\,
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7\,
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15\,
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23\,
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.counter_cry_7\,
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.counter_cry_15\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.counter_cry_23\,
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_11_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_11_21_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_11_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_11_23_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_12_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_12_22_0_\
        );

    \IN_MUX_bfv_17_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_3_0_\
        );

    \IN_MUX_bfv_17_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_17_4_0_\
        );

    \IN_MUX_bfv_17_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_17_5_0_\
        );

    \IN_MUX_bfv_17_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_17_6_0_\
        );

    \IN_MUX_bfv_17_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_7_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_17_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_15\,
            carryinitout => \bfn_17_21_0_\
        );

    \IN_MUX_bfv_17_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_23\,
            carryinitout => \bfn_17_22_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_15_12_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_17_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_23_0_\
        );

    \IN_MUX_bfv_17_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryinitout => \bfn_17_24_0_\
        );

    \IN_MUX_bfv_17_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryinitout => \bfn_17_25_0_\
        );

    \IN_MUX_bfv_17_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryinitout => \bfn_17_26_0_\
        );

    \IN_MUX_bfv_12_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_23_0_\
        );

    \IN_MUX_bfv_12_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            carryinitout => \bfn_12_24_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            carryinitout => \bfn_15_24_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21626\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21641\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__29003\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst1.stoper_tr.un2_start_0_g\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__24539\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_tr.un2_start_0_g\
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__49010\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_163_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__42106\,
            CLKHFEN => \N__42110\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__42218\,
            RGB2PWM => \N__23027\,
            RGB1 => rgb_g_wire,
            CURREN => \N__42779\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__23327\,
            RGB0PWM => \N__53465\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_0_c_inv_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21794\,
            in2 => \_gnd_net_\,
            in3 => \N__21809\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_1_c_inv_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21938\,
            in2 => \_gnd_net_\,
            in3 => \N__21953\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_2_c_inv_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21932\,
            in1 => \N__21917\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_3_c_inv_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21911\,
            in1 => \N__21896\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_4_c_inv_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21875\,
            in2 => \_gnd_net_\,
            in3 => \N__21890\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_5_c_inv_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21854\,
            in2 => \_gnd_net_\,
            in3 => \N__21869\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_6_c_inv_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21833\,
            in2 => \_gnd_net_\,
            in3 => \N__21848\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_7_c_inv_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21815\,
            in2 => \_gnd_net_\,
            in3 => \N__21827\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_8_c_inv_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22085\,
            in2 => \_gnd_net_\,
            in3 => \N__22097\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_9_c_inv_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22064\,
            in2 => \_gnd_net_\,
            in3 => \N__22079\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_10_c_inv_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22043\,
            in2 => \_gnd_net_\,
            in3 => \N__22058\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_10\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_11_c_inv_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22022\,
            in2 => \_gnd_net_\,
            in3 => \N__22037\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_12_c_inv_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22001\,
            in2 => \_gnd_net_\,
            in3 => \N__22016\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_12\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_13_c_inv_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21980\,
            in2 => \_gnd_net_\,
            in3 => \N__21995\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_13\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_14_c_inv_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21959\,
            in2 => \_gnd_net_\,
            in3 => \N__21974\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_15_c_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22172\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_16_c_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22133\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_16_c_RNIL8HR_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22223\,
            in2 => \_gnd_net_\,
            in3 => \N__22121\,
            lcout => \pwm_generator_inst.un22_threshold_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_17_c_RNINCJR_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22217\,
            in2 => \_gnd_net_\,
            in3 => \N__22118\,
            lcout => \pwm_generator_inst.un18_threshold1_18\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_18_c_RNIPGLR_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23507\,
            in2 => \_gnd_net_\,
            in3 => \N__22115\,
            lcout => \pwm_generator_inst.un18_threshold1_19\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_18\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_19_c_RNIRKNR_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22229\,
            in2 => \_gnd_net_\,
            in3 => \N__22112\,
            lcout => \pwm_generator_inst.un18_threshold1_20\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_19\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_20_c_RNIK7IS_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22205\,
            in2 => \_gnd_net_\,
            in3 => \N__22109\,
            lcout => \pwm_generator_inst.un18_threshold1_21\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_20\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_21_c_RNIMBKS_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22211\,
            in2 => \_gnd_net_\,
            in3 => \N__22106\,
            lcout => \pwm_generator_inst.un18_threshold1_22\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_21\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_22_c_RNIOFMS_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23186\,
            in2 => \_gnd_net_\,
            in3 => \N__22103\,
            lcout => \pwm_generator_inst.un18_threshold1_23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_22\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_23_c_RNIQJOS_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23141\,
            in2 => \_gnd_net_\,
            in3 => \N__22100\,
            lcout => \pwm_generator_inst.un18_threshold1_24\,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_24_c_RNISNQS_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23333\,
            in2 => \_gnd_net_\,
            in3 => \N__22235\,
            lcout => \pwm_generator_inst.un18_threshold1_25\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_24\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_25_c_RNIK5UE2_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010011010"
        )
    port map (
            in0 => \N__22556\,
            in1 => \N__23273\,
            in2 => \N__23899\,
            in3 => \N__22232\,
            lcout => \pwm_generator_inst.N_188_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_0_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23965\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_0_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23233\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_0_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23005\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_0_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23806\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_0_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23920\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_15_c_RNO_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22199\,
            in2 => \N__22187\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_15\,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_16_c_RNO_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22163\,
            in2 => \N__22151\,
            in3 => \N__22124\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_16\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22502\,
            in2 => \N__22490\,
            in3 => \N__22472\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22469\,
            in2 => \N__22457\,
            in3 => \N__22436\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22433\,
            in2 => \N__22421\,
            in3 => \N__22403\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRROZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22400\,
            in2 => \N__22388\,
            in3 => \N__22370\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22367\,
            in2 => \N__22352\,
            in3 => \N__22337\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22334\,
            in2 => \N__22319\,
            in3 => \N__22304\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22301\,
            in2 => \N__22286\,
            in3 => \N__22271\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0\,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22268\,
            in2 => \N__22253\,
            in3 => \N__22238\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22604\,
            in2 => \N__22589\,
            in3 => \N__22574\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPF_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23477\,
            in2 => \N__22571\,
            in3 => \N__22547\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_12_c_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22544\,
            in2 => \N__23492\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_13_c_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23481\,
            in2 => \N__22532\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_14_c_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22517\,
            in2 => \N__23493\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_15_c_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23485\,
            in2 => \N__23042\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJ1_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23357\,
            in2 => \_gnd_net_\,
            in3 => \N__22505\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29879\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_20_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CC_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22862\,
            in2 => \_gnd_net_\,
            in3 => \N__22829\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CCZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DC_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41989\,
            in2 => \N__22826\,
            in3 => \N__22790\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DCZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI77EC_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22787\,
            in2 => \N__42095\,
            in3 => \N__22754\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI77ECZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FC_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22751\,
            in2 => \_gnd_net_\,
            in3 => \N__22721\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FCZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGC_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22718\,
            in2 => \N__42096\,
            in3 => \N__22691\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGCZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHC_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22688\,
            in2 => \_gnd_net_\,
            in3 => \N__22655\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHCZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFIC_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22652\,
            in2 => \_gnd_net_\,
            in3 => \N__22622\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFICZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FO_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36773\,
            in3 => \N__22607\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FOZ0\,
            ltout => OPEN,
            carryin => \bfn_1_21_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDI8_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36722\,
            in3 => \N__22982\,
            lcout => \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDIZ0Z8\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_RNISHK8_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36665\,
            in3 => \N__22967\,
            lcout => \pwm_generator_inst.un3_threshold_cry_9_c_RNISHKZ0Z8\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_RNI59G7_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36608\,
            in3 => \N__22952\,
            lcout => \pwm_generator_inst.un3_threshold_cry_10_c_RNI59GZ0Z7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DI7_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37142\,
            in2 => \_gnd_net_\,
            in3 => \N__22937\,
            lcout => \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DIZ0Z7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HK7_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37106\,
            in2 => \_gnd_net_\,
            in3 => \N__22922\,
            lcout => \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HKZ0Z7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLM7_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37076\,
            in2 => \_gnd_net_\,
            in3 => \N__22907\,
            lcout => \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLMZ0Z7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPO7_LC_1_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37037\,
            in2 => \_gnd_net_\,
            in3 => \N__22892\,
            lcout => \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPOZ0Z7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQ7_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37001\,
            in2 => \_gnd_net_\,
            in3 => \N__22877\,
            lcout => \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQZ0Z7\,
            ltout => OPEN,
            carryin => \bfn_1_22_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1T7_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36968\,
            in2 => \_gnd_net_\,
            in3 => \N__23078\,
            lcout => \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1TZ0Z7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFD_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36932\,
            in2 => \_gnd_net_\,
            in3 => \N__23063\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFDZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJF_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37334\,
            in2 => \_gnd_net_\,
            in3 => \N__23060\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSON_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37316\,
            in1 => \N__23057\,
            in2 => \N__36896\,
            in3 => \N__23045\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSONZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNO_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__23494\,
            in1 => \N__23398\,
            in2 => \_gnd_net_\,
            in3 => \N__23380\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.N_112_i_i_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__26992\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53463\,
            lcout => \N_112_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNITBL3_9_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24048\,
            in1 => \N__24087\,
            in2 => \_gnd_net_\,
            in3 => \N__24222\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_2_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__23676\,
            in1 => \N__23631\,
            in2 => \N__23708\,
            in3 => \N__23135\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_6_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23021\,
            in1 => \N__24126\,
            in2 => \N__23015\,
            in3 => \N__24184\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_0_c_RNIIIGF3_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__23108\,
            in1 => \N__23889\,
            in2 => \N__23129\,
            in3 => \N__23012\,
            lcout => \pwm_generator_inst.N_180_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIRPD2_0_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23781\,
            in2 => \_gnd_net_\,
            in3 => \N__23754\,
            lcout => \pwm_generator_inst.un1_counterlto2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_0_c_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23245\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_0_THRU_LUT4_0_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42190\,
            in2 => \N__23125\,
            in3 => \N__23099\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_1_THRU_LUT4_0_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23536\,
            in2 => \N__42342\,
            in3 => \N__23096\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_2_THRU_LUT4_0_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42194\,
            in2 => \N__23998\,
            in3 => \N__23093\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_3_THRU_LUT4_0_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23938\,
            in2 => \N__42343\,
            in3 => \N__23090\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_4_THRU_LUT4_0_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42198\,
            in2 => \N__23830\,
            in3 => \N__23087\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_5_THRU_LUT4_0_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23206\,
            in2 => \N__42344\,
            in3 => \N__23084\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_6_THRU_LUT4_0_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42202\,
            in2 => \N__23177\,
            in3 => \N__23081\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_7_THRU_LUT4_0_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23263\,
            in2 => \N__42189\,
            in3 => \N__23279\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_16_0_\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_8_THRU_LUT4_0_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23276\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_7_c_RNI5Q6H3_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__23348\,
            in1 => \N__23885\,
            in2 => \N__23267\,
            in3 => \N__23252\,
            lcout => \pwm_generator_inst.N_187_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_16_c_RNI9O983_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23884\,
            in1 => \N__23246\,
            in2 => \_gnd_net_\,
            in3 => \N__23234\,
            lcout => \pwm_generator_inst.N_179_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_5_c_RNIT9UG3_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010101010"
        )
    port map (
            in0 => \N__23195\,
            in1 => \N__23222\,
            in2 => \N__23213\,
            in3 => \N__23879\,
            lcout => \pwm_generator_inst.N_185_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_0_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23194\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_6_c_RNI1I2H3_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010101010"
        )
    port map (
            in0 => \N__23150\,
            in1 => \N__23176\,
            in2 => \N__23162\,
            in3 => \N__23880\,
            lcout => \pwm_generator_inst.N_186_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_0_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23149\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_axb_16_1_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23495\,
            in2 => \_gnd_net_\,
            in3 => \N__23432\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un5_threshold_add_1_axb_16Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNICSGJ1_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010010110"
        )
    port map (
            in0 => \N__23417\,
            in1 => \N__23405\,
            in2 => \N__23387\,
            in3 => \N__23384\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_0_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23344\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.un8_start_stop_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__53464\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26996\,
            lcout => un8_start_stop,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23318\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23588\,
            in1 => \N__23785\,
            in2 => \_gnd_net_\,
            in3 => \N__23291\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_12_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__53843\,
            ce => 'H',
            sr => \N__53396\
        );

    \pwm_generator_inst.counter_1_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23582\,
            in1 => \N__23758\,
            in2 => \_gnd_net_\,
            in3 => \N__23288\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__53843\,
            ce => 'H',
            sr => \N__53396\
        );

    \pwm_generator_inst.counter_2_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23589\,
            in1 => \N__23706\,
            in2 => \_gnd_net_\,
            in3 => \N__23285\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__53843\,
            ce => 'H',
            sr => \N__53396\
        );

    \pwm_generator_inst.counter_3_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23583\,
            in1 => \N__23677\,
            in2 => \_gnd_net_\,
            in3 => \N__23282\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__53843\,
            ce => 'H',
            sr => \N__53396\
        );

    \pwm_generator_inst.counter_4_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23590\,
            in1 => \N__23632\,
            in2 => \_gnd_net_\,
            in3 => \N__23606\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__53843\,
            ce => 'H',
            sr => \N__53396\
        );

    \pwm_generator_inst.counter_5_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23584\,
            in1 => \N__24223\,
            in2 => \_gnd_net_\,
            in3 => \N__23603\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__53843\,
            ce => 'H',
            sr => \N__53396\
        );

    \pwm_generator_inst.counter_6_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23591\,
            in1 => \N__24183\,
            in2 => \_gnd_net_\,
            in3 => \N__23600\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__53843\,
            ce => 'H',
            sr => \N__53396\
        );

    \pwm_generator_inst.counter_7_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23585\,
            in1 => \N__24127\,
            in2 => \_gnd_net_\,
            in3 => \N__23597\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__53843\,
            ce => 'H',
            sr => \N__53396\
        );

    \pwm_generator_inst.counter_8_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23587\,
            in1 => \N__24091\,
            in2 => \_gnd_net_\,
            in3 => \N__23594\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_13_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__53837\,
            ce => 'H',
            sr => \N__53405\
        );

    \pwm_generator_inst.counter_9_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__24052\,
            in1 => \N__23586\,
            in2 => \_gnd_net_\,
            in3 => \N__23552\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53837\,
            ce => 'H',
            sr => \N__53405\
        );

    \pwm_generator_inst.un22_threshold_1_cry_1_c_RNIMQKF3_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010010111000"
        )
    port map (
            in0 => \N__23549\,
            in1 => \N__23900\,
            in2 => \N__23525\,
            in3 => \N__23543\,
            lcout => \pwm_generator_inst.N_181_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_0_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23521\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_2_c_RNIQ2PF3_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__24002\,
            in1 => \N__23981\,
            in2 => \N__23975\,
            in3 => \N__23902\,
            lcout => \pwm_generator_inst.N_182_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_3_c_RNILPLG3_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__23954\,
            in1 => \N__23903\,
            in2 => \N__23948\,
            in3 => \N__23927\,
            lcout => \pwm_generator_inst.N_183_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_4_c_RNIP1QG3_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__23909\,
            in1 => \N__23901\,
            in2 => \N__23837\,
            in3 => \N__23813\,
            lcout => \pwm_generator_inst.N_184_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23765\,
            in2 => \N__23795\,
            in3 => \N__23786\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_3_15_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23759\,
            in1 => \N__23723\,
            in2 => \N__23738\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23684\,
            in2 => \N__23717\,
            in3 => \N__23707\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23678\,
            in1 => \N__23648\,
            in2 => \N__23657\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23612\,
            in2 => \N__23642\,
            in3 => \N__23633\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24224\,
            in1 => \N__24191\,
            in2 => \N__24203\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24185\,
            in1 => \N__24149\,
            in2 => \N__24164\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24107\,
            in2 => \N__24143\,
            in3 => \N__24128\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24071\,
            in2 => \N__24101\,
            in3 => \N__24092\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_3_16_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24032\,
            in2 => \N__24065\,
            in3 => \N__24053\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24026\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53817\,
            ce => 'H',
            sr => \N__53415\
        );

    \CONSTANT_ONE_LUT4_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_15_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26351\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53824\,
            ce => \N__24456\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_12_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26120\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53818\,
            ce => \N__24448\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_14_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26372\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53819\,
            ce => \N__24443\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_28_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27793\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53809\,
            ce => \N__24447\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_2_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26045\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53801\,
            ce => \N__24457\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_13_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26393\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53801\,
            ce => \N__24457\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_25_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28499\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53794\,
            ce => \N__24455\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25866\,
            in2 => \_gnd_net_\,
            in3 => \N__24615\,
            lcout => \phase_controller_inst2.stoper_tr.un4_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101111111001100"
        )
    port map (
            in0 => \N__26820\,
            in1 => \N__24569\,
            in2 => \N__26797\,
            in3 => \N__24620\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53847\,
            ce => 'H',
            sr => \N__53344\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24621\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53847\,
            ce => 'H',
            sr => \N__53344\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__41094\,
            in1 => \N__41133\,
            in2 => \_gnd_net_\,
            in3 => \N__38558\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53844\,
            ce => 'H',
            sr => \N__53348\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__25874\,
            in1 => \N__53460\,
            in2 => \_gnd_net_\,
            in3 => \N__24623\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25875\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_4_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__26884\,
            in1 => \N__26910\,
            in2 => \_gnd_net_\,
            in3 => \N__26976\,
            lcout => \phase_controller_inst1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53830\,
            ce => 'H',
            sr => \N__53363\
        );

    \phase_controller_inst1.start_flag_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__26975\,
            in1 => \_gnd_net_\,
            in2 => \N__26917\,
            in3 => \N__26883\,
            lcout => \phase_controller_inst1.start_flagZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53830\,
            ce => 'H',
            sr => \N__53363\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__24511\,
            in1 => \N__24961\,
            in2 => \N__24322\,
            in3 => \N__24706\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__24512\,
            in1 => \N__24960\,
            in2 => \N__24323\,
            in3 => \N__24705\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010110010"
        )
    port map (
            in0 => \N__24233\,
            in1 => \N__24924\,
            in2 => \N__24484\,
            in3 => \N__24943\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010111011"
        )
    port map (
            in0 => \N__24232\,
            in1 => \N__24925\,
            in2 => \N__24485\,
            in3 => \N__24942\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_23_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30191\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53825\,
            ce => \N__24406\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__24524\,
            in1 => \N__24889\,
            in2 => \N__24269\,
            in3 => \N__24907\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__24523\,
            in1 => \N__24888\,
            in2 => \N__24268\,
            in3 => \N__24906\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001110"
        )
    port map (
            in0 => \N__24335\,
            in1 => \N__24497\,
            in2 => \N__24854\,
            in3 => \N__24871\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111010101111"
        )
    port map (
            in0 => \N__24334\,
            in1 => \N__24496\,
            in2 => \N__24853\,
            in3 => \N__24870\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33116\,
            in1 => \N__41053\,
            in2 => \_gnd_net_\,
            in3 => \N__31772\,
            lcout => \elapsed_time_ns_1_RNI0CQBB_0_31\,
            ltout => \elapsed_time_ns_1_RNI0CQBB_0_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_0_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__41020\,
            in1 => \_gnd_net_\,
            in2 => \N__24245\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53810\,
            ce => \N__24407\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32777\,
            in1 => \N__24242\,
            in2 => \_gnd_net_\,
            in3 => \N__31773\,
            lcout => \elapsed_time_ns_1_RNI1BOBB_0_14\,
            ltout => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24236\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26089\,
            in1 => \N__32963\,
            in2 => \_gnd_net_\,
            in3 => \N__31774\,
            lcout => \elapsed_time_ns_1_RNI1CPBB_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__24287\,
            in1 => \N__24785\,
            in2 => \N__24815\,
            in3 => \N__24278\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__24286\,
            in1 => \N__24784\,
            in2 => \N__24814\,
            in3 => \N__24277\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__24296\,
            in1 => \N__24731\,
            in2 => \N__24761\,
            in3 => \N__24305\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__24295\,
            in1 => \N__24730\,
            in2 => \N__24760\,
            in3 => \N__24304\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_19_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26267\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53802\,
            ce => \N__24437\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_1_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26060\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53795\,
            ce => \N__24439\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_11_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26138\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53795\,
            ce => \N__24439\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_7_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26203\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53795\,
            ce => \N__24439\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_18_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26288\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53795\,
            ce => \N__24439\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_16_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26330\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53795\,
            ce => \N__24439\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_17_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26309\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53795\,
            ce => \N__24439\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_27_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26420\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53795\,
            ce => \N__24439\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_3_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26027\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53795\,
            ce => \N__24439\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_4_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26008\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53788\,
            ce => \N__24438\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_5_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26236\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53788\,
            ce => \N__24438\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_6_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26218\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53788\,
            ce => \N__24438\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_21_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30224\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53788\,
            ce => \N__24438\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_8_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26186\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53788\,
            ce => \N__24438\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_10_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26153\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53788\,
            ce => \N__24438\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26059\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53786\,
            ce => \N__40956\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_11_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26134\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53786\,
            ce => \N__40956\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_12_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26113\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53786\,
            ce => \N__40956\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_13_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26386\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53786\,
            ce => \N__40956\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_14_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26365\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53786\,
            ce => \N__40956\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_15_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26344\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53786\,
            ce => \N__40956\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_2_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26041\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53786\,
            ce => \N__40956\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_3_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26026\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53786\,
            ce => \N__40956\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_4_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26012\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53783\,
            ce => \N__40955\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_5_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26240\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53783\,
            ce => \N__40955\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_6_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26222\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53783\,
            ce => \N__40955\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_7_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26204\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53783\,
            ce => \N__40955\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_8_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26185\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53783\,
            ce => \N__40955\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_9_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26167\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53783\,
            ce => \N__40955\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_10_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26152\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53783\,
            ce => \N__40955\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_24_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28510\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53782\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_20_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30238\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53782\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_26_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28465\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53782\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_9_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26171\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53782\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_22_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30205\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53782\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_16_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26329\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53778\,
            ce => \N__40954\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__28651\,
            in1 => \N__28640\,
            in2 => \N__28619\,
            in3 => \N__28585\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_17_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26308\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53778\,
            ce => \N__40954\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__26483\,
            in1 => \N__24557\,
            in2 => \N__26510\,
            in3 => \N__24548\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_18_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26284\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53778\,
            ce => \N__40954\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__26482\,
            in1 => \N__24556\,
            in2 => \N__26509\,
            in3 => \N__24547\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_19_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26263\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53778\,
            ce => \N__40954\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_27_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26416\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53766\,
            ce => \N__40937\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__24582\,
            in1 => \N__24622\,
            in2 => \_gnd_net_\,
            in3 => \N__25873\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__26576\,
            in1 => \N__26787\,
            in2 => \N__26600\,
            in3 => \N__26834\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53848\,
            ce => 'H',
            sr => \N__53339\
        );

    \phase_controller_inst2.state_3_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100011111111"
        )
    port map (
            in0 => \N__24652\,
            in1 => \N__26970\,
            in2 => \N__24640\,
            in3 => \N__26564\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53848\,
            ce => 'H',
            sr => \N__53339\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011100000"
        )
    port map (
            in0 => \N__26595\,
            in1 => \N__24583\,
            in2 => \N__24662\,
            in3 => \N__25828\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53848\,
            ce => 'H',
            sr => \N__53339\
        );

    \phase_controller_inst2.state_4_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010000010101010"
        )
    port map (
            in0 => \N__24653\,
            in1 => \_gnd_net_\,
            in2 => \N__24641\,
            in3 => \N__26971\,
            lcout => \phase_controller_inst2.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53848\,
            ce => 'H',
            sr => \N__53339\
        );

    \phase_controller_inst2.start_flag_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__26969\,
            in1 => \N__24651\,
            in2 => \_gnd_net_\,
            in3 => \N__24639\,
            lcout => \phase_controller_inst2.start_flagZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53848\,
            ce => 'H',
            sr => \N__53339\
        );

    \phase_controller_inst2.stoper_tr.running_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111001001110"
        )
    port map (
            in0 => \N__24619\,
            in1 => \N__24584\,
            in2 => \N__25876\,
            in3 => \N__25829\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53848\,
            ce => 'H',
            sr => \N__53339\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26723\,
            in2 => \_gnd_net_\,
            in3 => \N__26651\,
            lcout => \phase_controller_inst2.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26698\,
            in2 => \_gnd_net_\,
            in3 => \N__30675\,
            lcout => \phase_controller_inst2.stoper_hc.un4_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.counter_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25259\,
            in1 => \N__25135\,
            in2 => \N__25808\,
            in3 => \N__25807\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_0\,
            clk => \N__53838\,
            ce => \N__25157\,
            sr => \N__53345\
        );

    \phase_controller_inst2.stoper_tr.counter_1_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25267\,
            in1 => \N__25102\,
            in2 => \_gnd_net_\,
            in3 => \N__24563\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_1\,
            clk => \N__53838\,
            ce => \N__25157\,
            sr => \N__53345\
        );

    \phase_controller_inst2.stoper_tr.counter_2_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25260\,
            in1 => \N__25066\,
            in2 => \_gnd_net_\,
            in3 => \N__24560\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_2\,
            clk => \N__53838\,
            ce => \N__25157\,
            sr => \N__53345\
        );

    \phase_controller_inst2.stoper_tr.counter_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25268\,
            in1 => \N__25027\,
            in2 => \_gnd_net_\,
            in3 => \N__24689\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_3\,
            clk => \N__53838\,
            ce => \N__25157\,
            sr => \N__53345\
        );

    \phase_controller_inst2.stoper_tr.counter_4_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25261\,
            in1 => \N__24988\,
            in2 => \_gnd_net_\,
            in3 => \N__24686\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_4\,
            clk => \N__53838\,
            ce => \N__25157\,
            sr => \N__53345\
        );

    \phase_controller_inst2.stoper_tr.counter_5_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25269\,
            in1 => \N__25546\,
            in2 => \_gnd_net_\,
            in3 => \N__24683\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_5\,
            clk => \N__53838\,
            ce => \N__25157\,
            sr => \N__53345\
        );

    \phase_controller_inst2.stoper_tr.counter_6_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25262\,
            in1 => \N__25495\,
            in2 => \_gnd_net_\,
            in3 => \N__24680\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_6\,
            clk => \N__53838\,
            ce => \N__25157\,
            sr => \N__53345\
        );

    \phase_controller_inst2.stoper_tr.counter_7_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25270\,
            in1 => \N__25456\,
            in2 => \_gnd_net_\,
            in3 => \N__24677\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_7\,
            clk => \N__53838\,
            ce => \N__25157\,
            sr => \N__53345\
        );

    \phase_controller_inst2.stoper_tr.counter_8_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25258\,
            in1 => \N__25432\,
            in2 => \_gnd_net_\,
            in3 => \N__24674\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_8\,
            clk => \N__53831\,
            ce => \N__25158\,
            sr => \N__53349\
        );

    \phase_controller_inst2.stoper_tr.counter_9_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25274\,
            in1 => \N__25384\,
            in2 => \_gnd_net_\,
            in3 => \N__24671\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_9\,
            clk => \N__53831\,
            ce => \N__25158\,
            sr => \N__53349\
        );

    \phase_controller_inst2.stoper_tr.counter_10_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25255\,
            in1 => \N__25348\,
            in2 => \_gnd_net_\,
            in3 => \N__24668\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_10\,
            clk => \N__53831\,
            ce => \N__25158\,
            sr => \N__53349\
        );

    \phase_controller_inst2.stoper_tr.counter_11_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25271\,
            in1 => \N__25312\,
            in2 => \_gnd_net_\,
            in3 => \N__24665\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_11\,
            clk => \N__53831\,
            ce => \N__25158\,
            sr => \N__53349\
        );

    \phase_controller_inst2.stoper_tr.counter_12_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25256\,
            in1 => \N__25771\,
            in2 => \_gnd_net_\,
            in3 => \N__24827\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_12\,
            clk => \N__53831\,
            ce => \N__25158\,
            sr => \N__53349\
        );

    \phase_controller_inst2.stoper_tr.counter_13_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25272\,
            in1 => \N__25747\,
            in2 => \_gnd_net_\,
            in3 => \N__24824\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_13\,
            clk => \N__53831\,
            ce => \N__25158\,
            sr => \N__53349\
        );

    \phase_controller_inst2.stoper_tr.counter_14_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25257\,
            in1 => \N__25708\,
            in2 => \_gnd_net_\,
            in3 => \N__24821\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_14\,
            clk => \N__53831\,
            ce => \N__25158\,
            sr => \N__53349\
        );

    \phase_controller_inst2.stoper_tr.counter_15_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25273\,
            in1 => \N__25669\,
            in2 => \_gnd_net_\,
            in3 => \N__24818\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_15\,
            clk => \N__53831\,
            ce => \N__25158\,
            sr => \N__53349\
        );

    \phase_controller_inst2.stoper_tr.counter_16_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25283\,
            in1 => \N__24802\,
            in2 => \_gnd_net_\,
            in3 => \N__24788\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_16\,
            clk => \N__53826\,
            ce => \N__25159\,
            sr => \N__53357\
        );

    \phase_controller_inst2.stoper_tr.counter_17_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25263\,
            in1 => \N__24778\,
            in2 => \_gnd_net_\,
            in3 => \N__24764\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_17\,
            clk => \N__53826\,
            ce => \N__25159\,
            sr => \N__53357\
        );

    \phase_controller_inst2.stoper_tr.counter_18_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25284\,
            in1 => \N__24748\,
            in2 => \_gnd_net_\,
            in3 => \N__24734\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_18\,
            clk => \N__53826\,
            ce => \N__25159\,
            sr => \N__53357\
        );

    \phase_controller_inst2.stoper_tr.counter_19_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25264\,
            in1 => \N__24724\,
            in2 => \_gnd_net_\,
            in3 => \N__24710\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_19\,
            clk => \N__53826\,
            ce => \N__25159\,
            sr => \N__53357\
        );

    \phase_controller_inst2.stoper_tr.counter_20_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25285\,
            in1 => \N__24707\,
            in2 => \_gnd_net_\,
            in3 => \N__24692\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_20\,
            clk => \N__53826\,
            ce => \N__25159\,
            sr => \N__53357\
        );

    \phase_controller_inst2.stoper_tr.counter_21_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25265\,
            in1 => \N__24962\,
            in2 => \_gnd_net_\,
            in3 => \N__24947\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_21\,
            clk => \N__53826\,
            ce => \N__25159\,
            sr => \N__53357\
        );

    \phase_controller_inst2.stoper_tr.counter_22_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25286\,
            in1 => \N__24944\,
            in2 => \_gnd_net_\,
            in3 => \N__24929\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_22\,
            clk => \N__53826\,
            ce => \N__25159\,
            sr => \N__53357\
        );

    \phase_controller_inst2.stoper_tr.counter_23_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25266\,
            in1 => \N__24926\,
            in2 => \_gnd_net_\,
            in3 => \N__24911\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_23\,
            clk => \N__53826\,
            ce => \N__25159\,
            sr => \N__53357\
        );

    \phase_controller_inst2.stoper_tr.counter_24_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25275\,
            in1 => \N__24908\,
            in2 => \_gnd_net_\,
            in3 => \N__24893\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_24\,
            clk => \N__53820\,
            ce => \N__25160\,
            sr => \N__53364\
        );

    \phase_controller_inst2.stoper_tr.counter_25_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25279\,
            in1 => \N__24890\,
            in2 => \_gnd_net_\,
            in3 => \N__24875\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_25\,
            clk => \N__53820\,
            ce => \N__25160\,
            sr => \N__53364\
        );

    \phase_controller_inst2.stoper_tr.counter_26_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25276\,
            in1 => \N__24872\,
            in2 => \_gnd_net_\,
            in3 => \N__24857\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_26\,
            clk => \N__53820\,
            ce => \N__25160\,
            sr => \N__53364\
        );

    \phase_controller_inst2.stoper_tr.counter_27_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25280\,
            in1 => \N__24852\,
            in2 => \_gnd_net_\,
            in3 => \N__24833\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_27\,
            clk => \N__53820\,
            ce => \N__25160\,
            sr => \N__53364\
        );

    \phase_controller_inst2.stoper_tr.counter_28_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25277\,
            in1 => \N__25900\,
            in2 => \_gnd_net_\,
            in3 => \N__24830\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_28\,
            clk => \N__53820\,
            ce => \N__25160\,
            sr => \N__53364\
        );

    \phase_controller_inst2.stoper_tr.counter_29_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25281\,
            in1 => \N__25924\,
            in2 => \_gnd_net_\,
            in3 => \N__25292\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_29\,
            clk => \N__53820\,
            ce => \N__25160\,
            sr => \N__53364\
        );

    \phase_controller_inst2.stoper_tr.counter_30_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25278\,
            in1 => \N__34086\,
            in2 => \_gnd_net_\,
            in3 => \N__25289\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_29\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_30\,
            clk => \N__53820\,
            ce => \N__25160\,
            sr => \N__53364\
        );

    \phase_controller_inst2.stoper_tr.counter_31_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25282\,
            in1 => \N__34116\,
            in2 => \_gnd_net_\,
            in3 => \N__25163\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53820\,
            ce => \N__25160\,
            sr => \N__53364\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25142\,
            in2 => \N__25121\,
            in3 => \N__25136\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25112\,
            in2 => \N__25088\,
            in3 => \N__25103\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25079\,
            in2 => \N__25052\,
            in3 => \N__25067\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25040\,
            in2 => \N__25013\,
            in3 => \N__25028\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25004\,
            in2 => \N__24974\,
            in3 => \N__24992\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25547\,
            in1 => \N__25532\,
            in2 => \N__25520\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25511\,
            in2 => \N__25481\,
            in3 => \N__25499\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25469\,
            in2 => \N__25442\,
            in3 => \N__25460\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25433\,
            in1 => \N__25418\,
            in2 => \N__25406\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25397\,
            in2 => \N__25370\,
            in3 => \N__25385\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25361\,
            in2 => \N__25334\,
            in3 => \N__25349\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25298\,
            in2 => \N__25325\,
            in3 => \N__25313\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25784\,
            in2 => \N__25757\,
            in3 => \N__25772\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25748\,
            in1 => \N__25733\,
            in2 => \N__25721\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25709\,
            in1 => \N__25694\,
            in2 => \N__25682\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25673\,
            in1 => \N__25640\,
            in2 => \N__25655\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25634\,
            in2 => \N__25628\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25616\,
            in2 => \N__25610\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25598\,
            in2 => \N__25586\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25571\,
            in2 => \N__25562\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25994\,
            in2 => \N__25985\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25970\,
            in2 => \N__25961\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25886\,
            in2 => \N__25943\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34043\,
            in2 => \N__26075\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25946\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100000000"
        )
    port map (
            in0 => \N__25931\,
            in1 => \_gnd_net_\,
            in2 => \N__25910\,
            in3 => \N__34062\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__34061\,
            in1 => \N__25930\,
            in2 => \_gnd_net_\,
            in3 => \N__25906\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25880\,
            in2 => \_gnd_net_\,
            in3 => \N__25819\,
            lcout => \phase_controller_inst2.stoper_tr.counter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26099\,
            in1 => \N__32753\,
            in2 => \_gnd_net_\,
            in3 => \N__31787\,
            lcout => \elapsed_time_ns_1_RNI2COBB_0_15\,
            ltout => \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26093\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26090\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__34124\,
            in1 => \N__34097\,
            in2 => \_gnd_net_\,
            in3 => \N__34063\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26066\,
            in2 => \N__41016\,
            in3 => \N__41073\,
            lcout => \phase_controller_inst1.stoper_tr.measured_delay_tr_i_31\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27245\,
            in1 => \N__27241\,
            in2 => \N__42595\,
            in3 => \N__26048\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_1,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27221\,
            in1 => \N__27220\,
            in2 => \N__42599\,
            in3 => \N__26030\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_2,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27199\,
            in1 => \N__27200\,
            in2 => \N__42596\,
            in3 => \N__26015\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_3,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27170\,
            in1 => \N__27166\,
            in2 => \N__42600\,
            in3 => \N__25997\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_4,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27145\,
            in1 => \N__27146\,
            in2 => \N__42597\,
            in3 => \N__26225\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_5,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27125\,
            in1 => \N__27124\,
            in2 => \N__42601\,
            in3 => \N__26207\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_6,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27110\,
            in1 => \N__27109\,
            in2 => \N__42598\,
            in3 => \N__26189\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_7,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27095\,
            in1 => \N__27094\,
            in2 => \N__42362\,
            in3 => \N__26174\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_8,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27434\,
            in1 => \N__27430\,
            in2 => \N__42359\,
            in3 => \N__26156\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_9,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27410\,
            in1 => \N__27406\,
            in2 => \N__42363\,
            in3 => \N__26141\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_10,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27373\,
            in1 => \N__27374\,
            in2 => \N__42356\,
            in3 => \N__26123\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_11,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27344\,
            in1 => \N__27340\,
            in2 => \N__42360\,
            in3 => \N__26102\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_12,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27319\,
            in1 => \N__27320\,
            in2 => \N__42357\,
            in3 => \N__26375\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_13,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27299\,
            in1 => \N__27298\,
            in2 => \N__42361\,
            in3 => \N__26354\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_14,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27284\,
            in1 => \N__27283\,
            in2 => \N__42358\,
            in3 => \N__26333\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_15,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27268\,
            in1 => \N__27269\,
            in2 => \N__42452\,
            in3 => \N__26312\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_16,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27632\,
            in1 => \N__27628\,
            in2 => \N__42223\,
            in3 => \N__26291\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_17,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27599\,
            in1 => \N__27595\,
            in2 => \N__42453\,
            in3 => \N__26270\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_18,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27574\,
            in1 => \N__27575\,
            in2 => \N__42224\,
            in3 => \N__26249\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_19,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27548\,
            in1 => \N__27544\,
            in2 => \N__42454\,
            in3 => \N__26246\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_20,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27526\,
            in1 => \N__27527\,
            in2 => \N__42225\,
            in3 => \N__26243\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_21,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27506\,
            in1 => \N__27505\,
            in2 => \N__42455\,
            in3 => \N__26435\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_22,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27491\,
            in1 => \N__27490\,
            in2 => \N__42226\,
            in3 => \N__26432\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_23,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27476\,
            in1 => \N__27475\,
            in2 => \N__42219\,
            in3 => \N__26429\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_24,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27455\,
            in1 => \N__27451\,
            in2 => \N__42221\,
            in3 => \N__26426\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_25,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27851\,
            in1 => \N__27847\,
            in2 => \N__42220\,
            in3 => \N__26423\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_26,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27826\,
            in1 => \N__27827\,
            in2 => \N__42222\,
            in3 => \N__26402\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_27,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26399\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.counter_0_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28827\,
            in1 => \N__27757\,
            in2 => \N__28352\,
            in3 => \N__28351\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_0\,
            clk => \N__53774\,
            ce => \N__26627\,
            sr => \N__53413\
        );

    \phase_controller_inst1.stoper_tr.counter_1_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28831\,
            in1 => \N__27721\,
            in2 => \_gnd_net_\,
            in3 => \N__26396\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_1\,
            clk => \N__53774\,
            ce => \N__26627\,
            sr => \N__53413\
        );

    \phase_controller_inst1.stoper_tr.counter_2_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28828\,
            in1 => \N__27682\,
            in2 => \_gnd_net_\,
            in3 => \N__26462\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_2\,
            clk => \N__53774\,
            ce => \N__26627\,
            sr => \N__53413\
        );

    \phase_controller_inst1.stoper_tr.counter_3_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28832\,
            in1 => \N__27646\,
            in2 => \_gnd_net_\,
            in3 => \N__26459\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_3\,
            clk => \N__53774\,
            ce => \N__26627\,
            sr => \N__53413\
        );

    \phase_controller_inst1.stoper_tr.counter_4_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28829\,
            in1 => \N__28093\,
            in2 => \_gnd_net_\,
            in3 => \N__26456\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_4\,
            clk => \N__53774\,
            ce => \N__26627\,
            sr => \N__53413\
        );

    \phase_controller_inst1.stoper_tr.counter_5_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28833\,
            in1 => \N__28066\,
            in2 => \_gnd_net_\,
            in3 => \N__26453\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_5\,
            clk => \N__53774\,
            ce => \N__26627\,
            sr => \N__53413\
        );

    \phase_controller_inst1.stoper_tr.counter_6_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28830\,
            in1 => \N__28033\,
            in2 => \_gnd_net_\,
            in3 => \N__26450\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_6\,
            clk => \N__53774\,
            ce => \N__26627\,
            sr => \N__53413\
        );

    \phase_controller_inst1.stoper_tr.counter_7_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28834\,
            in1 => \N__27997\,
            in2 => \_gnd_net_\,
            in3 => \N__26447\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_7\,
            clk => \N__53774\,
            ce => \N__26627\,
            sr => \N__53413\
        );

    \phase_controller_inst1.stoper_tr.counter_8_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28813\,
            in1 => \N__27946\,
            in2 => \_gnd_net_\,
            in3 => \N__26444\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_21_0_\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_8\,
            clk => \N__53767\,
            ce => \N__26626\,
            sr => \N__53416\
        );

    \phase_controller_inst1.stoper_tr.counter_9_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28838\,
            in1 => \N__27913\,
            in2 => \_gnd_net_\,
            in3 => \N__26441\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_9\,
            clk => \N__53767\,
            ce => \N__26626\,
            sr => \N__53416\
        );

    \phase_controller_inst1.stoper_tr.counter_10_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28810\,
            in1 => \N__27874\,
            in2 => \_gnd_net_\,
            in3 => \N__26438\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_10\,
            clk => \N__53767\,
            ce => \N__26626\,
            sr => \N__53416\
        );

    \phase_controller_inst1.stoper_tr.counter_11_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28835\,
            in1 => \N__28315\,
            in2 => \_gnd_net_\,
            in3 => \N__26531\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_11\,
            clk => \N__53767\,
            ce => \N__26626\,
            sr => \N__53416\
        );

    \phase_controller_inst1.stoper_tr.counter_12_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28811\,
            in1 => \N__28276\,
            in2 => \_gnd_net_\,
            in3 => \N__26528\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_12\,
            clk => \N__53767\,
            ce => \N__26626\,
            sr => \N__53416\
        );

    \phase_controller_inst1.stoper_tr.counter_13_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28836\,
            in1 => \N__28255\,
            in2 => \_gnd_net_\,
            in3 => \N__26525\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_13\,
            clk => \N__53767\,
            ce => \N__26626\,
            sr => \N__53416\
        );

    \phase_controller_inst1.stoper_tr.counter_14_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28812\,
            in1 => \N__28219\,
            in2 => \_gnd_net_\,
            in3 => \N__26522\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_14\,
            clk => \N__53767\,
            ce => \N__26626\,
            sr => \N__53416\
        );

    \phase_controller_inst1.stoper_tr.counter_15_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28837\,
            in1 => \N__28183\,
            in2 => \_gnd_net_\,
            in3 => \N__26519\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_15\,
            clk => \N__53767\,
            ce => \N__26626\,
            sr => \N__53416\
        );

    \phase_controller_inst1.stoper_tr.counter_16_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28806\,
            in1 => \N__28614\,
            in2 => \_gnd_net_\,
            in3 => \N__26516\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_22_0_\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_16\,
            clk => \N__53763\,
            ce => \N__26625\,
            sr => \N__53417\
        );

    \phase_controller_inst1.stoper_tr.counter_17_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28814\,
            in1 => \N__28639\,
            in2 => \_gnd_net_\,
            in3 => \N__26513\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_17\,
            clk => \N__53763\,
            ce => \N__26625\,
            sr => \N__53417\
        );

    \phase_controller_inst1.stoper_tr.counter_18_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28807\,
            in1 => \N__26502\,
            in2 => \_gnd_net_\,
            in3 => \N__26486\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_18\,
            clk => \N__53763\,
            ce => \N__26625\,
            sr => \N__53417\
        );

    \phase_controller_inst1.stoper_tr.counter_19_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28815\,
            in1 => \N__26481\,
            in2 => \_gnd_net_\,
            in3 => \N__26465\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_19\,
            clk => \N__53763\,
            ce => \N__26625\,
            sr => \N__53417\
        );

    \phase_controller_inst1.stoper_tr.counter_20_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28808\,
            in1 => \N__30432\,
            in2 => \_gnd_net_\,
            in3 => \N__26558\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_20\,
            clk => \N__53763\,
            ce => \N__26625\,
            sr => \N__53417\
        );

    \phase_controller_inst1.stoper_tr.counter_21_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28816\,
            in1 => \N__30480\,
            in2 => \_gnd_net_\,
            in3 => \N__26555\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_21\,
            clk => \N__53763\,
            ce => \N__26625\,
            sr => \N__53417\
        );

    \phase_controller_inst1.stoper_tr.counter_22_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28809\,
            in1 => \N__30339\,
            in2 => \_gnd_net_\,
            in3 => \N__26552\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_22\,
            clk => \N__53763\,
            ce => \N__26625\,
            sr => \N__53417\
        );

    \phase_controller_inst1.stoper_tr.counter_23_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28817\,
            in1 => \N__30367\,
            in2 => \_gnd_net_\,
            in3 => \N__26549\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_23\,
            clk => \N__53763\,
            ce => \N__26625\,
            sr => \N__53417\
        );

    \phase_controller_inst1.stoper_tr.counter_24_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28780\,
            in1 => \N__28879\,
            in2 => \_gnd_net_\,
            in3 => \N__26546\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_23_0_\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_24\,
            clk => \N__53756\,
            ce => \N__26624\,
            sr => \N__53418\
        );

    \phase_controller_inst1.stoper_tr.counter_25_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28784\,
            in1 => \N__28912\,
            in2 => \_gnd_net_\,
            in3 => \N__26543\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_25\,
            clk => \N__53756\,
            ce => \N__26624\,
            sr => \N__53418\
        );

    \phase_controller_inst1.stoper_tr.counter_26_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28781\,
            in1 => \N__28409\,
            in2 => \_gnd_net_\,
            in3 => \N__26540\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_26\,
            clk => \N__53756\,
            ce => \N__26624\,
            sr => \N__53418\
        );

    \phase_controller_inst1.stoper_tr.counter_27_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28785\,
            in1 => \N__28451\,
            in2 => \_gnd_net_\,
            in3 => \N__26537\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_27\,
            clk => \N__53756\,
            ce => \N__26624\,
            sr => \N__53418\
        );

    \phase_controller_inst1.stoper_tr.counter_28_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28782\,
            in1 => \N__28561\,
            in2 => \_gnd_net_\,
            in3 => \N__26534\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_28\,
            clk => \N__53756\,
            ce => \N__26624\,
            sr => \N__53418\
        );

    \phase_controller_inst1.stoper_tr.counter_29_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28786\,
            in1 => \N__28545\,
            in2 => \_gnd_net_\,
            in3 => \N__26636\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_29\,
            clk => \N__53756\,
            ce => \N__26624\,
            sr => \N__53418\
        );

    \phase_controller_inst1.stoper_tr.counter_30_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28783\,
            in1 => \N__28988\,
            in2 => \_gnd_net_\,
            in3 => \N__26633\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_29\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_30\,
            clk => \N__53756\,
            ce => \N__26624\,
            sr => \N__53418\
        );

    \phase_controller_inst1.stoper_tr.counter_31_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28787\,
            in1 => \N__28943\,
            in2 => \_gnd_net_\,
            in3 => \N__26630\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53756\,
            ce => \N__26624\,
            sr => \N__53418\
        );

    \phase_controller_inst2.S2_LC_8_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26798\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53735\,
            ce => 'H',
            sr => \N__53423\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30684\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__30683\,
            in1 => \N__26678\,
            in2 => \_gnd_net_\,
            in3 => \N__26707\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__26708\,
            in1 => \N__53458\,
            in2 => \_gnd_net_\,
            in3 => \N__30682\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_RNO_0_3_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__26752\,
            in1 => \N__28691\,
            in2 => \N__26599\,
            in3 => \N__26575\,
            lcout => \phase_controller_inst2.state_ns_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__26705\,
            in1 => \N__26758\,
            in2 => \N__28699\,
            in3 => \N__26730\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53839\,
            ce => 'H',
            sr => \N__53340\
        );

    \phase_controller_inst2.state_1_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__26833\,
            in1 => \N__26786\,
            in2 => \N__26731\,
            in3 => \N__26654\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53839\,
            ce => 'H',
            sr => \N__53340\
        );

    \phase_controller_inst2.stoper_hc.running_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111001001110"
        )
    port map (
            in0 => \N__26704\,
            in1 => \N__26676\,
            in2 => \N__30685\,
            in3 => \N__31122\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53839\,
            ce => 'H',
            sr => \N__53340\
        );

    \phase_controller_inst2.state_2_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__26759\,
            in1 => \N__28695\,
            in2 => \N__26732\,
            in3 => \N__26653\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53839\,
            ce => 'H',
            sr => \N__53340\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26706\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53839\,
            ce => 'H',
            sr => \N__53340\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000000000"
        )
    port map (
            in0 => \N__26677\,
            in1 => \N__26652\,
            in2 => \N__31124\,
            in3 => \N__26660\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53839\,
            ce => 'H',
            sr => \N__53340\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33311\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53832\,
            ce => \N__37649\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_11_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33460\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53832\,
            ce => \N__37649\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_28_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27794\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53827\,
            ce => \N__40966\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34307\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53821\,
            ce => \N__34247\,
            sr => \N__53350\
        );

    \phase_controller_inst1.state_RNO_0_3_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__29592\,
            in1 => \N__49118\,
            in2 => \N__26867\,
            in3 => \N__26851\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.state_ns_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_3_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111110001111"
        )
    port map (
            in0 => \N__26980\,
            in1 => \N__26918\,
            in2 => \N__26894\,
            in3 => \N__26891\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53811\,
            ce => 'H',
            sr => \N__53358\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37249\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37276\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.un4_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__29019\,
            in1 => \N__26866\,
            in2 => \N__26870\,
            in3 => \N__28369\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53811\,
            ce => 'H',
            sr => \N__53358\
        );

    \phase_controller_inst1.state_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__26865\,
            in1 => \N__29614\,
            in2 => \N__30731\,
            in3 => \N__26852\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53811\,
            ce => 'H',
            sr => \N__53358\
        );

    \phase_controller_inst1.start_timer_tr_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101011111010"
        )
    port map (
            in0 => \N__29756\,
            in1 => \N__29613\,
            in2 => \N__37287\,
            in3 => \N__30729\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53811\,
            ce => 'H',
            sr => \N__53358\
        );

    \phase_controller_inst1.stoper_tr.running_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001001110010"
        )
    port map (
            in0 => \N__37277\,
            in1 => \N__37250\,
            in2 => \N__29026\,
            in3 => \N__28370\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53811\,
            ce => 'H',
            sr => \N__53358\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29785\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32552\,
            in1 => \N__26843\,
            in2 => \_gnd_net_\,
            in3 => \N__31734\,
            lcout => \elapsed_time_ns_1_RNIJI91B_0_7\,
            ltout => \elapsed_time_ns_1_RNIJI91B_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26837\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32638\,
            in1 => \N__27064\,
            in2 => \N__32621\,
            in3 => \N__27073\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34340\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53796\,
            ce => \N__34246\,
            sr => \N__53368\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31732\,
            in1 => \N__27044\,
            in2 => \_gnd_net_\,
            in3 => \N__27074\,
            lcout => \elapsed_time_ns_1_RNIDC91B_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31733\,
            in1 => \N__27023\,
            in2 => \_gnd_net_\,
            in3 => \N__27065\,
            lcout => \elapsed_time_ns_1_RNIED91B_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31727\,
            in1 => \N__27053\,
            in2 => \_gnd_net_\,
            in3 => \N__32639\,
            lcout => \elapsed_time_ns_1_RNIFE91B_0_3\,
            ltout => \elapsed_time_ns_1_RNIFE91B_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27047\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27043\,
            in1 => \N__41072\,
            in2 => \N__27032\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27011\,
            in2 => \_gnd_net_\,
            in3 => \N__27022\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27005\,
            in2 => \_gnd_net_\,
            in3 => \N__26999\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29966\,
            in2 => \_gnd_net_\,
            in3 => \N__27224\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29891\,
            in2 => \_gnd_net_\,
            in3 => \N__27203\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29807\,
            in2 => \_gnd_net_\,
            in3 => \N__27182\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27179\,
            in2 => \_gnd_net_\,
            in3 => \N__27149\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29723\,
            in2 => \_gnd_net_\,
            in3 => \N__27128\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29792\,
            in2 => \_gnd_net_\,
            in3 => \N__27113\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30029\,
            in2 => \_gnd_net_\,
            in3 => \N__27098\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29948\,
            in2 => \_gnd_net_\,
            in3 => \N__27077\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30044\,
            in2 => \_gnd_net_\,
            in3 => \N__27413\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29741\,
            in2 => \_gnd_net_\,
            in3 => \N__27389\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27386\,
            in2 => \_gnd_net_\,
            in3 => \N__27356\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27353\,
            in3 => \N__27323\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30062\,
            in2 => \_gnd_net_\,
            in3 => \N__27302\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30014\,
            in3 => \N__27287\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30119\,
            in2 => \_gnd_net_\,
            in3 => \N__27272\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30401\,
            in2 => \_gnd_net_\,
            in3 => \N__27248\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29933\,
            in3 => \N__27611\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27608\,
            in2 => \_gnd_net_\,
            in3 => \N__27578\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31628\,
            in2 => \_gnd_net_\,
            in3 => \N__27557\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27554\,
            in2 => \_gnd_net_\,
            in3 => \N__27530\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29906\,
            in2 => \_gnd_net_\,
            in3 => \N__27509\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30077\,
            in2 => \_gnd_net_\,
            in3 => \N__27494\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0\,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30134\,
            in2 => \_gnd_net_\,
            in3 => \N__27479\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30092\,
            in2 => \_gnd_net_\,
            in3 => \N__27458\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30245\,
            in2 => \_gnd_net_\,
            in3 => \N__27854\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27767\,
            in2 => \_gnd_net_\,
            in3 => \N__27830\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29990\,
            in2 => \_gnd_net_\,
            in3 => \N__27809\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__27806\,
            in1 => \N__41074\,
            in2 => \_gnd_net_\,
            in3 => \N__27797\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30112\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27761\,
            in1 => \N__40985\,
            in2 => \N__27743\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27734\,
            in2 => \N__27707\,
            in3 => \N__27722\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27695\,
            in2 => \N__27668\,
            in3 => \N__27683\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27659\,
            in2 => \N__28112\,
            in3 => \N__27647\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28103\,
            in2 => \N__28079\,
            in3 => \N__28094\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28067\,
            in1 => \N__28052\,
            in2 => \N__28043\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28034\,
            in1 => \N__28019\,
            in2 => \N__28010\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28001\,
            in1 => \N__27983\,
            in2 => \N__27974\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27932\,
            in2 => \N__27965\,
            in3 => \N__27950\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27926\,
            in2 => \N__27899\,
            in3 => \N__27914\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27860\,
            in2 => \N__27890\,
            in3 => \N__27875\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28328\,
            in2 => \N__28301\,
            in3 => \N__28316\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28262\,
            in2 => \N__28292\,
            in3 => \N__28277\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28256\,
            in1 => \N__28241\,
            in2 => \N__28229\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28220\,
            in1 => \N__28205\,
            in2 => \N__28193\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28184\,
            in1 => \N__28169\,
            in2 => \N__28157\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28574\,
            in2 => \N__28148\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28133\,
            in2 => \N__28124\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30416\,
            in2 => \N__30170\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28523\,
            in2 => \N__30302\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28382\,
            in2 => \N__28853\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28478\,
            in2 => \N__28394\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28529\,
            in2 => \N__28337\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29039\,
            in2 => \N__28928\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28373\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37242\,
            in2 => \_gnd_net_\,
            in3 => \N__28363\,
            lcout => \phase_controller_inst1.stoper_tr.counter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__28567\,
            in1 => \N__28967\,
            in2 => \_gnd_net_\,
            in3 => \N__28546\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__28658\,
            in1 => \N__28638\,
            in2 => \N__28618\,
            in3 => \N__28592\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__28568\,
            in1 => \N__28968\,
            in2 => \_gnd_net_\,
            in3 => \N__28547\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__30385\,
            in1 => \N__30363\,
            in2 => \N__30343\,
            in3 => \N__30316\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_24_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28517\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53757\,
            ce => \N__40915\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_25_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28498\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53757\,
            ce => \N__40915\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011010100"
        )
    port map (
            in0 => \N__28450\,
            in1 => \N__28436\,
            in2 => \N__28424\,
            in3 => \N__28408\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_26_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28469\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53757\,
            ce => \N__40915\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011011101"
        )
    port map (
            in0 => \N__28449\,
            in1 => \N__28435\,
            in2 => \N__28423\,
            in3 => \N__28407\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__28861\,
            in1 => \N__28878\,
            in2 => \N__28916\,
            in3 => \N__28891\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__28941\,
            in1 => \N__28986\,
            in2 => \_gnd_net_\,
            in3 => \N__28972\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__29030\,
            in1 => \N__37293\,
            in2 => \_gnd_net_\,
            in3 => \N__37238\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__28987\,
            in1 => \_gnd_net_\,
            in2 => \N__28973\,
            in3 => \N__28942\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__28908\,
            in1 => \N__28892\,
            in2 => \N__28880\,
            in3 => \N__28862\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37243\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S1_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28706\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53729\,
            ce => 'H',
            sr => \N__53424\
        );

    \phase_controller_inst2.stoper_hc.counter_0_LC_10_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29348\,
            in1 => \N__30619\,
            in2 => \N__30638\,
            in3 => \N__30637\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_2_0_\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_0\,
            clk => \N__53851\,
            ce => \N__29260\,
            sr => \N__53319\
        );

    \phase_controller_inst2.stoper_hc.counter_1_LC_10_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29390\,
            in1 => \N__30598\,
            in2 => \_gnd_net_\,
            in3 => \N__28661\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_1\,
            clk => \N__53851\,
            ce => \N__29260\,
            sr => \N__53319\
        );

    \phase_controller_inst2.stoper_hc.counter_2_LC_10_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29349\,
            in1 => \N__30571\,
            in2 => \_gnd_net_\,
            in3 => \N__29066\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_2\,
            clk => \N__53851\,
            ce => \N__29260\,
            sr => \N__53319\
        );

    \phase_controller_inst2.stoper_hc.counter_3_LC_10_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29391\,
            in1 => \N__30547\,
            in2 => \_gnd_net_\,
            in3 => \N__29063\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_3\,
            clk => \N__53851\,
            ce => \N__29260\,
            sr => \N__53319\
        );

    \phase_controller_inst2.stoper_hc.counter_4_LC_10_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29350\,
            in1 => \N__30526\,
            in2 => \_gnd_net_\,
            in3 => \N__29060\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_4\,
            clk => \N__53851\,
            ce => \N__29260\,
            sr => \N__53319\
        );

    \phase_controller_inst2.stoper_hc.counter_5_LC_10_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29392\,
            in1 => \N__30925\,
            in2 => \_gnd_net_\,
            in3 => \N__29057\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_5\,
            clk => \N__53851\,
            ce => \N__29260\,
            sr => \N__53319\
        );

    \phase_controller_inst2.stoper_hc.counter_6_LC_10_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29351\,
            in1 => \N__30904\,
            in2 => \_gnd_net_\,
            in3 => \N__29054\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_6\,
            clk => \N__53851\,
            ce => \N__29260\,
            sr => \N__53319\
        );

    \phase_controller_inst2.stoper_hc.counter_7_LC_10_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29393\,
            in1 => \N__30883\,
            in2 => \_gnd_net_\,
            in3 => \N__29051\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_7\,
            clk => \N__53851\,
            ce => \N__29260\,
            sr => \N__53319\
        );

    \phase_controller_inst2.stoper_hc.counter_8_LC_10_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29347\,
            in1 => \N__30859\,
            in2 => \_gnd_net_\,
            in3 => \N__29048\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_10_3_0_\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_8\,
            clk => \N__53849\,
            ce => \N__29256\,
            sr => \N__53321\
        );

    \phase_controller_inst2.stoper_hc.counter_9_LC_10_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29359\,
            in1 => \N__30835\,
            in2 => \_gnd_net_\,
            in3 => \N__29045\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_9\,
            clk => \N__53849\,
            ce => \N__29256\,
            sr => \N__53321\
        );

    \phase_controller_inst2.stoper_hc.counter_10_LC_10_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29344\,
            in1 => \N__30811\,
            in2 => \_gnd_net_\,
            in3 => \N__29042\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_10\,
            clk => \N__53849\,
            ce => \N__29256\,
            sr => \N__53321\
        );

    \phase_controller_inst2.stoper_hc.counter_11_LC_10_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29356\,
            in1 => \N__30787\,
            in2 => \_gnd_net_\,
            in3 => \N__29093\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_11\,
            clk => \N__53849\,
            ce => \N__29256\,
            sr => \N__53321\
        );

    \phase_controller_inst2.stoper_hc.counter_12_LC_10_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29345\,
            in1 => \N__30760\,
            in2 => \_gnd_net_\,
            in3 => \N__29090\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_12\,
            clk => \N__53849\,
            ce => \N__29256\,
            sr => \N__53321\
        );

    \phase_controller_inst2.stoper_hc.counter_13_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29357\,
            in1 => \N__31096\,
            in2 => \_gnd_net_\,
            in3 => \N__29087\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_13\,
            clk => \N__53849\,
            ce => \N__29256\,
            sr => \N__53321\
        );

    \phase_controller_inst2.stoper_hc.counter_14_LC_10_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29346\,
            in1 => \N__31069\,
            in2 => \_gnd_net_\,
            in3 => \N__29084\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_14\,
            clk => \N__53849\,
            ce => \N__29256\,
            sr => \N__53321\
        );

    \phase_controller_inst2.stoper_hc.counter_15_LC_10_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29358\,
            in1 => \N__31045\,
            in2 => \_gnd_net_\,
            in3 => \N__29081\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_15\,
            clk => \N__53849\,
            ce => \N__29256\,
            sr => \N__53321\
        );

    \phase_controller_inst2.stoper_hc.counter_16_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29352\,
            in1 => \N__29682\,
            in2 => \_gnd_net_\,
            in3 => \N__29078\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_10_4_0_\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_16\,
            clk => \N__53845\,
            ce => \N__29261\,
            sr => \N__53323\
        );

    \phase_controller_inst2.stoper_hc.counter_17_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29386\,
            in1 => \N__29715\,
            in2 => \_gnd_net_\,
            in3 => \N__29075\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_17\,
            clk => \N__53845\,
            ce => \N__29261\,
            sr => \N__53323\
        );

    \phase_controller_inst2.stoper_hc.counter_18_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29353\,
            in1 => \N__29490\,
            in2 => \_gnd_net_\,
            in3 => \N__29072\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_18\,
            clk => \N__53845\,
            ce => \N__29261\,
            sr => \N__53323\
        );

    \phase_controller_inst2.stoper_hc.counter_19_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29387\,
            in1 => \N__29463\,
            in2 => \_gnd_net_\,
            in3 => \N__29069\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_19\,
            clk => \N__53845\,
            ce => \N__29261\,
            sr => \N__53323\
        );

    \phase_controller_inst2.stoper_hc.counter_20_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29354\,
            in1 => \N__29136\,
            in2 => \_gnd_net_\,
            in3 => \N__29120\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_20\,
            clk => \N__53845\,
            ce => \N__29261\,
            sr => \N__53323\
        );

    \phase_controller_inst2.stoper_hc.counter_21_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29388\,
            in1 => \N__29160\,
            in2 => \_gnd_net_\,
            in3 => \N__29117\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_21\,
            clk => \N__53845\,
            ce => \N__29261\,
            sr => \N__53323\
        );

    \phase_controller_inst2.stoper_hc.counter_22_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29355\,
            in1 => \N__29439\,
            in2 => \_gnd_net_\,
            in3 => \N__29114\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_22\,
            clk => \N__53845\,
            ce => \N__29261\,
            sr => \N__53323\
        );

    \phase_controller_inst2.stoper_hc.counter_23_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29389\,
            in1 => \N__29415\,
            in2 => \_gnd_net_\,
            in3 => \N__29111\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_23\,
            clk => \N__53845\,
            ce => \N__29261\,
            sr => \N__53323\
        );

    \phase_controller_inst2.stoper_hc.counter_24_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29378\,
            in1 => \N__29547\,
            in2 => \_gnd_net_\,
            in3 => \N__29108\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_10_5_0_\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_24\,
            clk => \N__53840\,
            ce => \N__29249\,
            sr => \N__53326\
        );

    \phase_controller_inst2.stoper_hc.counter_25_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29383\,
            in1 => \N__29565\,
            in2 => \_gnd_net_\,
            in3 => \N__29105\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_25\,
            clk => \N__53840\,
            ce => \N__29249\,
            sr => \N__53326\
        );

    \phase_controller_inst2.stoper_hc.counter_26_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29379\,
            in1 => \N__29511\,
            in2 => \_gnd_net_\,
            in3 => \N__29102\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_26\,
            clk => \N__53840\,
            ce => \N__29249\,
            sr => \N__53326\
        );

    \phase_controller_inst2.stoper_hc.counter_27_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29384\,
            in1 => \N__29529\,
            in2 => \_gnd_net_\,
            in3 => \N__29099\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_27\,
            clk => \N__53840\,
            ce => \N__29249\,
            sr => \N__53326\
        );

    \phase_controller_inst2.stoper_hc.counter_28_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29380\,
            in1 => \N__29225\,
            in2 => \_gnd_net_\,
            in3 => \N__29096\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_28\,
            clk => \N__53840\,
            ce => \N__29249\,
            sr => \N__53326\
        );

    \phase_controller_inst2.stoper_hc.counter_29_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29385\,
            in1 => \N__29210\,
            in2 => \_gnd_net_\,
            in3 => \N__29399\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_29\,
            clk => \N__53840\,
            ce => \N__29249\,
            sr => \N__53326\
        );

    \phase_controller_inst2.stoper_hc.counter_30_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29381\,
            in1 => \N__29195\,
            in2 => \_gnd_net_\,
            in3 => \N__29396\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_29\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_30\,
            clk => \N__53840\,
            ce => \N__29249\,
            sr => \N__53326\
        );

    \phase_controller_inst2.stoper_hc.counter_31_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__29180\,
            in1 => \N__29382\,
            in2 => \_gnd_net_\,
            in3 => \N__29264\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53840\,
            ce => \N__29249\,
            sr => \N__53326\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__29224\,
            in1 => \N__29209\,
            in2 => \_gnd_net_\,
            in3 => \N__29649\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100101011"
        )
    port map (
            in0 => \N__33226\,
            in1 => \N__29161\,
            in2 => \N__29143\,
            in3 => \N__31219\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__29223\,
            in1 => \N__29208\,
            in2 => \_gnd_net_\,
            in3 => \N__29648\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__29650\,
            in1 => \N__29179\,
            in2 => \_gnd_net_\,
            in3 => \N__29193\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__29194\,
            in1 => \N__29178\,
            in2 => \_gnd_net_\,
            in3 => \N__29651\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101100100010"
        )
    port map (
            in0 => \N__33227\,
            in1 => \N__29162\,
            in2 => \N__29144\,
            in3 => \N__31220\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__29666\,
            in1 => \N__29467\,
            in2 => \N__29495\,
            in3 => \N__31238\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__31307\,
            in1 => \N__29567\,
            in2 => \N__31208\,
            in3 => \N__29549\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__31306\,
            in1 => \N__29566\,
            in2 => \N__31207\,
            in3 => \N__29548\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__29630\,
            in1 => \N__29531\,
            in2 => \N__31190\,
            in3 => \N__29513\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__29629\,
            in1 => \N__29530\,
            in2 => \N__31189\,
            in3 => \N__29512\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__29665\,
            in1 => \N__29491\,
            in2 => \N__29471\,
            in3 => \N__31234\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000100"
        )
    port map (
            in0 => \N__29441\,
            in1 => \N__31247\,
            in2 => \N__29423\,
            in3 => \N__31256\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100001101"
        )
    port map (
            in0 => \N__29440\,
            in1 => \N__31246\,
            in2 => \N__29422\,
            in3 => \N__31255\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__29717\,
            in1 => \N__29699\,
            in2 => \N__29690\,
            in3 => \N__31316\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_16_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33982\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53812\,
            ce => \N__33374\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__29716\,
            in1 => \N__29698\,
            in2 => \N__29689\,
            in3 => \N__31315\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_18_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34642\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53812\,
            ce => \N__33374\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_28_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36482\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53803\,
            ce => \N__33375\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_26_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33686\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53803\,
            ce => \N__33375\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_1_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__29773\,
            in1 => \N__29618\,
            in2 => \N__34154\,
            in3 => \N__30722\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53797\,
            ce => 'H',
            sr => \N__53346\
        );

    \phase_controller_inst1.state_2_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__29594\,
            in1 => \N__29774\,
            in2 => \N__49129\,
            in3 => \N__34153\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53797\,
            ce => 'H',
            sr => \N__53346\
        );

    \phase_controller_inst1.start_timer_hc_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__29593\,
            in1 => \N__34022\,
            in2 => \N__49128\,
            in3 => \N__29772\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53797\,
            ce => 'H',
            sr => \N__53346\
        );

    \phase_controller_inst1.stoper_hc.running_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111001001110"
        )
    port map (
            in0 => \N__34021\,
            in1 => \N__34198\,
            in2 => \N__34547\,
            in3 => \N__34178\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53797\,
            ce => 'H',
            sr => \N__53346\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34023\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53797\,
            ce => 'H',
            sr => \N__53346\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31759\,
            in1 => \N__30004\,
            in2 => \_gnd_net_\,
            in3 => \N__33143\,
            lcout => \elapsed_time_ns_1_RNIVAQBB_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31757\,
            in1 => \N__33011\,
            in2 => \_gnd_net_\,
            in3 => \N__29786\,
            lcout => \elapsed_time_ns_1_RNIV9PBB_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29920\,
            in1 => \N__32936\,
            in2 => \_gnd_net_\,
            in3 => \N__31758\,
            lcout => \elapsed_time_ns_1_RNI2DPBB_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29771\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34144\,
            lcout => \phase_controller_inst1.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29750\,
            in1 => \N__32804\,
            in2 => \_gnd_net_\,
            in3 => \N__31756\,
            lcout => \elapsed_time_ns_1_RNI0AOBB_0_13\,
            ltout => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29744\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__34197\,
            in1 => \N__34017\,
            in2 => \_gnd_net_\,
            in3 => \N__34527\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32527\,
            in1 => \N__29732\,
            in2 => \_gnd_net_\,
            in3 => \N__31735\,
            lcout => \elapsed_time_ns_1_RNIKJ91B_0_8\,
            ltout => \elapsed_time_ns_1_RNIKJ91B_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29726\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_i_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29878\,
            lcout => \pwm_generator_inst.un3_threshold_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31736\,
            in1 => \N__29960\,
            in2 => \_gnd_net_\,
            in3 => \N__32849\,
            lcout => \elapsed_time_ns_1_RNIU7OBB_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__32548\,
            in1 => \N__29828\,
            in2 => \N__32528\,
            in3 => \N__30158\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__33112\,
            in1 => \N__30143\,
            in2 => \N__29822\,
            in3 => \N__30284\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29816\,
            in2 => \N__29819\,
            in3 => \N__32573\,
            lcout => \elapsed_time_ns_1_RNIIH91B_0_6\,
            ltout => \elapsed_time_ns_1_RNIIH91B_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29810\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31729\,
            in1 => \N__29801\,
            in2 => \_gnd_net_\,
            in3 => \N__32507\,
            lcout => \elapsed_time_ns_1_RNILK91B_0_9\,
            ltout => \elapsed_time_ns_1_RNILK91B_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29795\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31730\,
            in1 => \N__30056\,
            in2 => \_gnd_net_\,
            in3 => \N__32825\,
            lcout => \elapsed_time_ns_1_RNIV8OBB_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32617\,
            in1 => \N__29975\,
            in2 => \_gnd_net_\,
            in3 => \N__31728\,
            lcout => \elapsed_time_ns_1_RNIGF91B_0_4\,
            ltout => \elapsed_time_ns_1_RNIGF91B_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29969\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29959\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31731\,
            in1 => \N__29942\,
            in2 => \_gnd_net_\,
            in3 => \N__33035\,
            lcout => \elapsed_time_ns_1_RNIU8PBB_0_20\,
            ltout => \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29936\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29921\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29900\,
            in1 => \N__32594\,
            in2 => \_gnd_net_\,
            in3 => \N__31766\,
            lcout => \elapsed_time_ns_1_RNIHG91B_0_5\,
            ltout => \elapsed_time_ns_1_RNIHG91B_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29894\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29885\,
            in1 => \N__32729\,
            in2 => \_gnd_net_\,
            in3 => \N__31768\,
            lcout => \elapsed_time_ns_1_RNI3DOBB_0_16\,
            ltout => \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30065\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30055\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31767\,
            in1 => \N__30038\,
            in2 => \_gnd_net_\,
            in3 => \N__32870\,
            lcout => \elapsed_time_ns_1_RNIT6OBB_0_10\,
            ltout => \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30032\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30023\,
            in1 => \N__32705\,
            in2 => \_gnd_net_\,
            in3 => \N__31769\,
            lcout => \elapsed_time_ns_1_RNI4EOBB_0_17\,
            ltout => \elapsed_time_ns_1_RNI4EOBB_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30017\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30005\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31771\,
            in1 => \N__29984\,
            in2 => \_gnd_net_\,
            in3 => \N__32891\,
            lcout => \elapsed_time_ns_1_RNI4FPBB_0_26\,
            ltout => \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29978\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31770\,
            in1 => \N__30128\,
            in2 => \_gnd_net_\,
            in3 => \N__33068\,
            lcout => \elapsed_time_ns_1_RNI5FOBB_0_18\,
            ltout => \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30122\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30113\,
            in1 => \N__33164\,
            in2 => \_gnd_net_\,
            in3 => \N__31781\,
            lcout => \elapsed_time_ns_1_RNI7IPBB_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31779\,
            in1 => \N__30101\,
            in2 => \_gnd_net_\,
            in3 => \N__33209\,
            lcout => \elapsed_time_ns_1_RNI5GPBB_0_27\,
            ltout => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30095\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30086\,
            in1 => \N__31778\,
            in2 => \_gnd_net_\,
            in3 => \N__32912\,
            lcout => \elapsed_time_ns_1_RNI3EPBB_0_25\,
            ltout => \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30080\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30071\,
            in1 => \N__33188\,
            in2 => \_gnd_net_\,
            in3 => \N__31780\,
            lcout => \elapsed_time_ns_1_RNI6HPBB_0_28\,
            ltout => \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30248\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_20_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30239\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53768\,
            ce => \N__40941\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_21_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30223\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53768\,
            ce => \N__40941\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_22_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30206\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53768\,
            ce => \N__40941\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_23_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30184\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53768\,
            ce => \N__40941\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__30487\,
            in1 => \N__30457\,
            in2 => \N__30443\,
            in3 => \N__30499\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32566\,
            in2 => \_gnd_net_\,
            in3 => \N__32587\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32839\,
            in1 => \N__32863\,
            in2 => \N__32503\,
            in3 => \N__32818\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32767\,
            in2 => \N__30146\,
            in3 => \N__32791\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010110010"
        )
    port map (
            in0 => \N__30503\,
            in1 => \N__30488\,
            in2 => \N__30461\,
            in3 => \N__30442\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30410\,
            in1 => \N__33047\,
            in2 => \_gnd_net_\,
            in3 => \N__31786\,
            lcout => \elapsed_time_ns_1_RNI6GOBB_0_19\,
            ltout => \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30404\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__30386\,
            in1 => \N__30371\,
            in2 => \N__30347\,
            in3 => \N__30317\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32698\,
            in1 => \N__32743\,
            in2 => \N__32725\,
            in3 => \N__33061\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33001\,
            in1 => \N__33025\,
            in2 => \N__32983\,
            in3 => \N__33046\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30293\,
            in1 => \N__30737\,
            in2 => \N__30287\,
            in3 => \N__30254\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_er_RNO_0_31_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30272\,
            in2 => \_gnd_net_\,
            in3 => \N__35980\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33202\,
            in1 => \N__32884\,
            in2 => \N__33184\,
            in3 => \N__32905\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33157\,
            in1 => \N__32950\,
            in2 => \N__32932\,
            in3 => \N__33133\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30730\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53727\,
            ce => 'H',
            sr => \N__53422\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30686\,
            in2 => \_gnd_net_\,
            in3 => \N__31123\,
            lcout => \phase_controller_inst2.stoper_hc.counter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30605\,
            in2 => \N__33404\,
            in3 => \N__30623\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_11_4_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33083\,
            in2 => \N__30584\,
            in3 => \N__30599\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33089\,
            in2 => \N__30557\,
            in3 => \N__30575\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30533\,
            in2 => \N__33242\,
            in3 => \N__30548\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30527\,
            in1 => \N__33266\,
            in2 => \N__30512\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30926\,
            in1 => \N__30911\,
            in2 => \N__33077\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30890\,
            in2 => \N__33251\,
            in3 => \N__30905\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30884\,
            in1 => \N__30869\,
            in2 => \N__33260\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30863\,
            in1 => \N__33410\,
            in2 => \N__30845\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30821\,
            in2 => \N__33275\,
            in3 => \N__30836\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33233\,
            in2 => \N__30797\,
            in3 => \N__30815\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33281\,
            in2 => \N__30773\,
            in3 => \N__30788\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30761\,
            in1 => \N__33215\,
            in2 => \N__30746\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31097\,
            in1 => \N__33416\,
            in2 => \N__31082\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33422\,
            in2 => \N__31055\,
            in3 => \N__31070\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31046\,
            in1 => \N__31031\,
            in2 => \N__33389\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31025\,
            in2 => \N__31013\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30998\,
            in2 => \N__30992\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30977\,
            in2 => \N__30971\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30962\,
            in2 => \N__30953\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30941\,
            in2 => \N__30935\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31172\,
            in2 => \N__31166\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31157\,
            in2 => \N__31151\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31142\,
            in2 => \N__31136\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31127\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_15_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33586\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53813\,
            ce => \N__37647\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_8_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33496\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53813\,
            ce => \N__37647\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_5_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33520\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53813\,
            ce => \N__37647\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_9_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33478\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53813\,
            ce => \N__37647\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_12_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33436\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53813\,
            ce => \N__37647\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_14_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33604\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53813\,
            ce => \N__37647\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_13_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33622\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53813\,
            ce => \N__37647\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_23_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33719\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53813\,
            ce => \N__37647\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_23_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33718\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53804\,
            ce => \N__33380\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_22_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33733\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53804\,
            ce => \N__33380\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_19_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33844\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53804\,
            ce => \N__33380\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_20_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33559\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53804\,
            ce => \N__33380\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_25_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33755\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53804\,
            ce => \N__33380\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_27_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33668\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53804\,
            ce => \N__33380\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_17_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34669\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53804\,
            ce => \N__33380\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_24_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33704\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53804\,
            ce => \N__33380\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__32180\,
            in1 => \N__31295\,
            in2 => \N__32210\,
            in3 => \N__31286\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_20_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33560\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53798\,
            ce => \N__37635\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__32179\,
            in1 => \N__31294\,
            in2 => \N__32209\,
            in3 => \N__31285\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_21_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33541\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53798\,
            ce => \N__37635\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__31277\,
            in1 => \N__32453\,
            in2 => \N__32483\,
            in3 => \N__31268\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_22_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33734\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53798\,
            ce => \N__37635\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__31276\,
            in1 => \N__32452\,
            in2 => \N__32482\,
            in3 => \N__31267\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__31382\,
            in1 => \N__32399\,
            in2 => \N__32428\,
            in3 => \N__33743\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_24_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33703\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53789\,
            ce => \N__37642\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__31381\,
            in1 => \N__32398\,
            in2 => \N__32429\,
            in3 => \N__33742\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__32348\,
            in1 => \N__31373\,
            in2 => \N__32375\,
            in3 => \N__31364\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_26_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33685\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53789\,
            ce => \N__37642\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__32347\,
            in1 => \N__31372\,
            in2 => \N__32374\,
            in3 => \N__31363\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_27_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33667\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53789\,
            ce => \N__37642\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37658\,
            in2 => \N__31355\,
            in3 => \N__31964\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31331\,
            in2 => \N__31346\,
            in3 => \N__31946\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33881\,
            in2 => \N__31325\,
            in3 => \N__31925\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33815\,
            in2 => \N__31487\,
            in3 => \N__31904\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33632\,
            in2 => \N__31475\,
            in3 => \N__31883\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32153\,
            in1 => \N__31463\,
            in2 => \N__31451\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31439\,
            in2 => \N__33857\,
            in3 => \N__32135\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32114\,
            in1 => \N__31433\,
            in2 => \N__33791\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32096\,
            in1 => \N__31427\,
            in2 => \N__31418\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31409\,
            in2 => \N__31400\,
            in3 => \N__32078\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33764\,
            in2 => \N__31391\,
            in3 => \N__32060\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31598\,
            in2 => \N__31616\,
            in3 => \N__32039\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31592\,
            in2 => \N__31580\,
            in3 => \N__32021\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31571\,
            in2 => \N__31562\,
            in3 => \N__32279\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32258\,
            in1 => \N__31550\,
            in2 => \N__31538\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32240\,
            in1 => \N__31514\,
            in2 => \N__31526\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33989\,
            in2 => \N__33908\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34649\,
            in2 => \N__34556\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31508\,
            in2 => \N__31499\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31862\,
            in2 => \N__31850\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31835\,
            in2 => \N__31826\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31814\,
            in2 => \N__31802\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31985\,
            in2 => \N__32000\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31991\,
            in2 => \N__36383\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31790\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31637\,
            in1 => \N__32987\,
            in2 => \_gnd_net_\,
            in3 => \N__31785\,
            lcout => \elapsed_time_ns_1_RNI0BPBB_0_22\,
            ltout => \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31631\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__32303\,
            in1 => \N__36405\,
            in2 => \_gnd_net_\,
            in3 => \N__32326\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__36407\,
            in1 => \N__36460\,
            in2 => \_gnd_net_\,
            in3 => \N__36430\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__32302\,
            in1 => \N__36406\,
            in2 => \_gnd_net_\,
            in3 => \N__32327\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34543\,
            in2 => \_gnd_net_\,
            in3 => \N__34167\,
            lcout => \phase_controller_inst1.stoper_hc.counter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.counter_0_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34493\,
            in1 => \N__31960\,
            in2 => \N__31979\,
            in3 => \N__31978\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_0\,
            clk => \N__53775\,
            ce => \N__32676\,
            sr => \N__53369\
        );

    \phase_controller_inst1.stoper_hc.counter_1_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34406\,
            in1 => \N__31942\,
            in2 => \_gnd_net_\,
            in3 => \N__31928\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_1\,
            clk => \N__53775\,
            ce => \N__32676\,
            sr => \N__53369\
        );

    \phase_controller_inst1.stoper_hc.counter_2_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34494\,
            in1 => \N__31921\,
            in2 => \_gnd_net_\,
            in3 => \N__31907\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_2\,
            clk => \N__53775\,
            ce => \N__32676\,
            sr => \N__53369\
        );

    \phase_controller_inst1.stoper_hc.counter_3_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34407\,
            in1 => \N__31903\,
            in2 => \_gnd_net_\,
            in3 => \N__31886\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_3\,
            clk => \N__53775\,
            ce => \N__32676\,
            sr => \N__53369\
        );

    \phase_controller_inst1.stoper_hc.counter_4_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34495\,
            in1 => \N__31879\,
            in2 => \_gnd_net_\,
            in3 => \N__31865\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_4\,
            clk => \N__53775\,
            ce => \N__32676\,
            sr => \N__53369\
        );

    \phase_controller_inst1.stoper_hc.counter_5_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34408\,
            in1 => \N__32152\,
            in2 => \_gnd_net_\,
            in3 => \N__32138\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_5\,
            clk => \N__53775\,
            ce => \N__32676\,
            sr => \N__53369\
        );

    \phase_controller_inst1.stoper_hc.counter_6_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34496\,
            in1 => \N__32131\,
            in2 => \_gnd_net_\,
            in3 => \N__32117\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_6\,
            clk => \N__53775\,
            ce => \N__32676\,
            sr => \N__53369\
        );

    \phase_controller_inst1.stoper_hc.counter_7_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34409\,
            in1 => \N__32113\,
            in2 => \_gnd_net_\,
            in3 => \N__32099\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_7\,
            clk => \N__53775\,
            ce => \N__32676\,
            sr => \N__53369\
        );

    \phase_controller_inst1.stoper_hc.counter_8_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34436\,
            in1 => \N__32095\,
            in2 => \_gnd_net_\,
            in3 => \N__32081\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_8\,
            clk => \N__53769\,
            ce => \N__32678\,
            sr => \N__53373\
        );

    \phase_controller_inst1.stoper_hc.counter_9_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34492\,
            in1 => \N__32077\,
            in2 => \_gnd_net_\,
            in3 => \N__32063\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_9\,
            clk => \N__53769\,
            ce => \N__32678\,
            sr => \N__53373\
        );

    \phase_controller_inst1.stoper_hc.counter_10_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34433\,
            in1 => \N__32056\,
            in2 => \_gnd_net_\,
            in3 => \N__32042\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_10\,
            clk => \N__53769\,
            ce => \N__32678\,
            sr => \N__53373\
        );

    \phase_controller_inst1.stoper_hc.counter_11_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34489\,
            in1 => \N__32038\,
            in2 => \_gnd_net_\,
            in3 => \N__32024\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_11\,
            clk => \N__53769\,
            ce => \N__32678\,
            sr => \N__53373\
        );

    \phase_controller_inst1.stoper_hc.counter_12_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34434\,
            in1 => \N__32017\,
            in2 => \_gnd_net_\,
            in3 => \N__32003\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_12\,
            clk => \N__53769\,
            ce => \N__32678\,
            sr => \N__53373\
        );

    \phase_controller_inst1.stoper_hc.counter_13_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34490\,
            in1 => \N__32275\,
            in2 => \_gnd_net_\,
            in3 => \N__32261\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_13\,
            clk => \N__53769\,
            ce => \N__32678\,
            sr => \N__53373\
        );

    \phase_controller_inst1.stoper_hc.counter_14_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34435\,
            in1 => \N__32257\,
            in2 => \_gnd_net_\,
            in3 => \N__32243\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_14\,
            clk => \N__53769\,
            ce => \N__32678\,
            sr => \N__53373\
        );

    \phase_controller_inst1.stoper_hc.counter_15_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34491\,
            in1 => \N__32239\,
            in2 => \_gnd_net_\,
            in3 => \N__32225\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_15\,
            clk => \N__53769\,
            ce => \N__32678\,
            sr => \N__53373\
        );

    \phase_controller_inst1.stoper_hc.counter_16_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34481\,
            in1 => \N__33922\,
            in2 => \_gnd_net_\,
            in3 => \N__32222\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_16\,
            clk => \N__53764\,
            ce => \N__32677\,
            sr => \N__53378\
        );

    \phase_controller_inst1.stoper_hc.counter_17_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34485\,
            in1 => \N__33949\,
            in2 => \_gnd_net_\,
            in3 => \N__32219\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_17\,
            clk => \N__53764\,
            ce => \N__32677\,
            sr => \N__53378\
        );

    \phase_controller_inst1.stoper_hc.counter_18_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34482\,
            in1 => \N__34570\,
            in2 => \_gnd_net_\,
            in3 => \N__32216\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_18\,
            clk => \N__53764\,
            ce => \N__32677\,
            sr => \N__53378\
        );

    \phase_controller_inst1.stoper_hc.counter_19_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34486\,
            in1 => \N__34591\,
            in2 => \_gnd_net_\,
            in3 => \N__32213\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_19\,
            clk => \N__53764\,
            ce => \N__32677\,
            sr => \N__53378\
        );

    \phase_controller_inst1.stoper_hc.counter_20_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34483\,
            in1 => \N__32197\,
            in2 => \_gnd_net_\,
            in3 => \N__32183\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_20\,
            clk => \N__53764\,
            ce => \N__32677\,
            sr => \N__53378\
        );

    \phase_controller_inst1.stoper_hc.counter_21_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34487\,
            in1 => \N__32170\,
            in2 => \_gnd_net_\,
            in3 => \N__32156\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_21\,
            clk => \N__53764\,
            ce => \N__32677\,
            sr => \N__53378\
        );

    \phase_controller_inst1.stoper_hc.counter_22_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34484\,
            in1 => \N__32470\,
            in2 => \_gnd_net_\,
            in3 => \N__32456\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_22\,
            clk => \N__53764\,
            ce => \N__32677\,
            sr => \N__53378\
        );

    \phase_controller_inst1.stoper_hc.counter_23_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34488\,
            in1 => \N__32446\,
            in2 => \_gnd_net_\,
            in3 => \N__32432\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_23\,
            clk => \N__53764\,
            ce => \N__32677\,
            sr => \N__53378\
        );

    \phase_controller_inst1.stoper_hc.counter_24_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34455\,
            in1 => \N__32416\,
            in2 => \_gnd_net_\,
            in3 => \N__32402\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_24\,
            clk => \N__53758\,
            ce => \N__32675\,
            sr => \N__53384\
        );

    \phase_controller_inst1.stoper_hc.counter_25_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34460\,
            in1 => \N__32392\,
            in2 => \_gnd_net_\,
            in3 => \N__32378\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_25\,
            clk => \N__53758\,
            ce => \N__32675\,
            sr => \N__53384\
        );

    \phase_controller_inst1.stoper_hc.counter_26_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34456\,
            in1 => \N__32367\,
            in2 => \_gnd_net_\,
            in3 => \N__32351\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_26\,
            clk => \N__53758\,
            ce => \N__32675\,
            sr => \N__53384\
        );

    \phase_controller_inst1.stoper_hc.counter_27_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34461\,
            in1 => \N__32346\,
            in2 => \_gnd_net_\,
            in3 => \N__32330\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_27\,
            clk => \N__53758\,
            ce => \N__32675\,
            sr => \N__53384\
        );

    \phase_controller_inst1.stoper_hc.counter_28_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34457\,
            in1 => \N__32320\,
            in2 => \_gnd_net_\,
            in3 => \N__32306\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_28\,
            clk => \N__53758\,
            ce => \N__32675\,
            sr => \N__53384\
        );

    \phase_controller_inst1.stoper_hc.counter_29_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34462\,
            in1 => \N__32296\,
            in2 => \_gnd_net_\,
            in3 => \N__32282\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_29\,
            clk => \N__53758\,
            ce => \N__32675\,
            sr => \N__53384\
        );

    \phase_controller_inst1.stoper_hc.counter_30_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34458\,
            in1 => \N__36429\,
            in2 => \_gnd_net_\,
            in3 => \N__32684\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_29\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_30\,
            clk => \N__53758\,
            ce => \N__32675\,
            sr => \N__53384\
        );

    \phase_controller_inst1.stoper_hc.counter_31_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__36456\,
            in1 => \N__34459\,
            in2 => \_gnd_net_\,
            in3 => \N__32681\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53758\,
            ce => \N__32675\,
            sr => \N__53384\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34881\,
            in2 => \N__34333\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_11_20_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__53752\,
            ce => \N__34259\,
            sr => \N__53390\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34860\,
            in2 => \N__34297\,
            in3 => \N__32597\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__53752\,
            ce => \N__34259\,
            sr => \N__53390\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34882\,
            in2 => \N__34840\,
            in3 => \N__32576\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__53752\,
            ce => \N__34259\,
            sr => \N__53390\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34812\,
            in2 => \N__34865\,
            in3 => \N__32555\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__53752\,
            ce => \N__34259\,
            sr => \N__53390\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34788\,
            in2 => \N__34841\,
            in3 => \N__32531\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__53752\,
            ce => \N__34259\,
            sr => \N__53390\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34764\,
            in2 => \N__34817\,
            in3 => \N__32510\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__53752\,
            ce => \N__34259\,
            sr => \N__53390\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34740\,
            in2 => \N__34793\,
            in3 => \N__32486\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__53752\,
            ce => \N__34259\,
            sr => \N__53390\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34716\,
            in2 => \N__34769\,
            in3 => \N__32852\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__53752\,
            ce => \N__34259\,
            sr => \N__53390\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34692\,
            in2 => \N__34745\,
            in3 => \N__32828\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_11_21_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__53747\,
            ce => \N__34269\,
            sr => \N__53400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35070\,
            in2 => \N__34721\,
            in3 => \N__32807\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__53747\,
            ce => \N__34269\,
            sr => \N__53400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35046\,
            in2 => \N__34697\,
            in3 => \N__32780\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__53747\,
            ce => \N__34269\,
            sr => \N__53400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35022\,
            in2 => \N__35075\,
            in3 => \N__32756\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__53747\,
            ce => \N__34269\,
            sr => \N__53400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34998\,
            in2 => \N__35051\,
            in3 => \N__32732\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__53747\,
            ce => \N__34269\,
            sr => \N__53400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34974\,
            in2 => \N__35027\,
            in3 => \N__32708\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__53747\,
            ce => \N__34269\,
            sr => \N__53400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34950\,
            in2 => \N__35003\,
            in3 => \N__32687\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__53747\,
            ce => \N__34269\,
            sr => \N__53400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34926\,
            in2 => \N__34979\,
            in3 => \N__33050\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__53747\,
            ce => \N__34269\,
            sr => \N__53400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34902\,
            in2 => \N__34955\,
            in3 => \N__33038\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__53742\,
            ce => \N__34271\,
            sr => \N__53406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35256\,
            in2 => \N__34931\,
            in3 => \N__33014\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__53742\,
            ce => \N__34271\,
            sr => \N__53406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35232\,
            in2 => \N__34907\,
            in3 => \N__32990\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__53742\,
            ce => \N__34271\,
            sr => \N__53406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35208\,
            in2 => \N__35261\,
            in3 => \N__32966\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__53742\,
            ce => \N__34271\,
            sr => \N__53406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35184\,
            in2 => \N__35237\,
            in3 => \N__32939\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__53742\,
            ce => \N__34271\,
            sr => \N__53406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35160\,
            in2 => \N__35213\,
            in3 => \N__32915\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__53742\,
            ce => \N__34271\,
            sr => \N__53406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35136\,
            in2 => \N__35189\,
            in3 => \N__32894\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__53742\,
            ce => \N__34271\,
            sr => \N__53406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35112\,
            in2 => \N__35165\,
            in3 => \N__32873\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__53742\,
            ce => \N__34271\,
            sr => \N__53406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35091\,
            in2 => \N__35141\,
            in3 => \N__33191\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_11_23_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__53737\,
            ce => \N__34270\,
            sr => \N__53410\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35661\,
            in2 => \N__35117\,
            in3 => \N__33167\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__53737\,
            ce => \N__34270\,
            sr => \N__53410\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35092\,
            in2 => \N__35642\,
            in3 => \N__33146\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__53737\,
            ce => \N__34270\,
            sr => \N__53410\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35494\,
            in2 => \N__35666\,
            in3 => \N__33122\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__53737\,
            ce => \N__34270\,
            sr => \N__53410\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33119\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53737\,
            ce => \N__34270\,
            sr => \N__53410\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_2_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33895\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53833\,
            ce => \N__33367\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_1_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33307\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53833\,
            ce => \N__33367\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_5_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33524\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53833\,
            ce => \N__33367\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_11_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33461\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53828\,
            ce => \N__33352\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_9_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33482\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53828\,
            ce => \N__33352\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_4_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33649\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53828\,
            ce => \N__33352\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_7_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33808\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53828\,
            ce => \N__33352\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_6_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33874\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53828\,
            ce => \N__33352\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_3_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33829\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53828\,
            ce => \N__33352\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_10_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33781\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53822\,
            ce => \N__33376\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_21_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33545\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53822\,
            ce => \N__33376\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_12_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33440\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53822\,
            ce => \N__33376\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_14_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33608\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53822\,
            ce => \N__33376\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_13_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33626\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53822\,
            ce => \N__33376\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_8_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33500\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53822\,
            ce => \N__33376\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_0_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37735\,
            in2 => \_gnd_net_\,
            in3 => \N__37680\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53822\,
            ce => \N__33376\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_15_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33590\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53822\,
            ce => \N__33376\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33317\,
            in2 => \N__37681\,
            in3 => \N__37719\,
            lcout => \phase_controller_inst1.stoper_hc.measured_delay_hc_i_31\,
            ltout => OPEN,
            carryin => \bfn_12_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36086\,
            in1 => \N__36085\,
            in2 => \N__42772\,
            in3 => \N__33290\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_1,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36065\,
            in1 => \N__36064\,
            in2 => \N__42776\,
            in3 => \N__33287\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_2,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36050\,
            in1 => \N__36049\,
            in2 => \N__42773\,
            in3 => \N__33284\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_3,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36035\,
            in1 => \N__36034\,
            in2 => \N__42777\,
            in3 => \N__33527\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_4,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36020\,
            in1 => \N__36019\,
            in2 => \N__42774\,
            in3 => \N__33509\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_5,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36005\,
            in1 => \N__36004\,
            in2 => \N__42778\,
            in3 => \N__33506\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_6,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36239\,
            in1 => \N__36238\,
            in2 => \N__42775\,
            in3 => \N__33503\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_7,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36224\,
            in1 => \N__36223\,
            in2 => \N__42770\,
            in3 => \N__33485\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_8,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36209\,
            in1 => \N__36208\,
            in2 => \N__42767\,
            in3 => \N__33467\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_9,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36194\,
            in1 => \N__36193\,
            in2 => \N__42771\,
            in3 => \N__33464\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_10,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36179\,
            in1 => \N__36178\,
            in2 => \N__42764\,
            in3 => \N__33443\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_11,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36155\,
            in1 => \N__36154\,
            in2 => \N__42768\,
            in3 => \N__33425\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_12,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36140\,
            in1 => \N__36139\,
            in2 => \N__42765\,
            in3 => \N__33611\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_13,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36125\,
            in1 => \N__36124\,
            in2 => \N__42769\,
            in3 => \N__33593\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_14,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36110\,
            in1 => \N__36109\,
            in2 => \N__42766\,
            in3 => \N__33575\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_15,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36368\,
            in1 => \N__36367\,
            in2 => \N__42705\,
            in3 => \N__33572\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_16,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36353\,
            in1 => \N__36352\,
            in2 => \N__42709\,
            in3 => \N__33569\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_17,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36338\,
            in1 => \N__36337\,
            in2 => \N__42706\,
            in3 => \N__33566\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_18,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36314\,
            in1 => \N__36313\,
            in2 => \N__42710\,
            in3 => \N__33563\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_19,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36299\,
            in1 => \N__36298\,
            in2 => \N__42707\,
            in3 => \N__33548\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_20,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36284\,
            in1 => \N__36283\,
            in2 => \N__42711\,
            in3 => \N__33530\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_21,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36269\,
            in1 => \N__36268\,
            in2 => \N__42708\,
            in3 => \N__33722\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_22,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36254\,
            in1 => \N__36253\,
            in2 => \N__42712\,
            in3 => \N__33707\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_23,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36557\,
            in1 => \N__36556\,
            in2 => \N__42630\,
            in3 => \N__33692\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_24,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36542\,
            in1 => \N__36541\,
            in2 => \N__42632\,
            in3 => \N__33689\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_25,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36527\,
            in1 => \N__36526\,
            in2 => \N__42631\,
            in3 => \N__33671\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_26,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36512\,
            in1 => \N__36511\,
            in2 => \N__42633\,
            in3 => \N__33656\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_27,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33653\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_4_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33650\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53787\,
            ce => \N__37622\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_2_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33899\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53787\,
            ce => \N__37622\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_6_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33875\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53787\,
            ce => \N__37622\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_19_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33848\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53787\,
            ce => \N__37622\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_3_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33833\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53787\,
            ce => \N__37622\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_7_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33809\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53787\,
            ce => \N__37622\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_10_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33782\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53787\,
            ce => \N__37622\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_25_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33754\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53787\,
            ce => \N__37622\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__34359\,
            in1 => \_gnd_net_\,
            in2 => \N__48854\,
            in3 => \N__48877\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_168_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__48878\,
            in1 => \N__34360\,
            in2 => \_gnd_net_\,
            in3 => \N__48853\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53784\,
            ce => 'H',
            sr => \N__53341\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34358\,
            in2 => \_gnd_net_\,
            in3 => \N__48849\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_167_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34030\,
            in2 => \_gnd_net_\,
            in3 => \N__34546\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un4_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__34205\,
            in1 => \N__34143\,
            in2 => \N__34181\,
            in3 => \N__34174\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53784\,
            ce => 'H',
            sr => \N__53341\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__34123\,
            in1 => \N__34093\,
            in2 => \_gnd_net_\,
            in3 => \N__34070\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__34031\,
            in1 => \N__53459\,
            in2 => \_gnd_net_\,
            in3 => \N__34545\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49943\,
            in1 => \N__39049\,
            in2 => \N__49756\,
            in3 => \N__39011\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__33965\,
            in1 => \N__33956\,
            in2 => \N__33935\,
            in3 => \N__34658\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_16_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33983\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53779\,
            ce => \N__37600\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__33964\,
            in1 => \N__33955\,
            in2 => \N__33934\,
            in3 => \N__34657\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_17_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34673\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53779\,
            ce => \N__37600\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__34625\,
            in1 => \N__34616\,
            in2 => \N__34603\,
            in3 => \N__34577\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_18_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34643\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53779\,
            ce => \N__37600\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__34624\,
            in1 => \N__34615\,
            in2 => \N__34604\,
            in3 => \N__34576\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34544\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34361\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35586\,
            in1 => \N__34326\,
            in2 => \_gnd_net_\,
            in3 => \N__34310\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__53751\,
            ce => \N__35458\,
            sr => \N__53379\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35621\,
            in1 => \N__34290\,
            in2 => \_gnd_net_\,
            in3 => \N__34274\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__53751\,
            ce => \N__35458\,
            sr => \N__53379\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35587\,
            in1 => \N__34883\,
            in2 => \_gnd_net_\,
            in3 => \N__34868\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__53751\,
            ce => \N__35458\,
            sr => \N__53379\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35622\,
            in1 => \N__34861\,
            in2 => \_gnd_net_\,
            in3 => \N__34844\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__53751\,
            ce => \N__35458\,
            sr => \N__53379\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35588\,
            in1 => \N__34839\,
            in2 => \_gnd_net_\,
            in3 => \N__34820\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__53751\,
            ce => \N__35458\,
            sr => \N__53379\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35623\,
            in1 => \N__34813\,
            in2 => \_gnd_net_\,
            in3 => \N__34796\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__53751\,
            ce => \N__35458\,
            sr => \N__53379\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35589\,
            in1 => \N__34789\,
            in2 => \_gnd_net_\,
            in3 => \N__34772\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__53751\,
            ce => \N__35458\,
            sr => \N__53379\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35624\,
            in1 => \N__34765\,
            in2 => \_gnd_net_\,
            in3 => \N__34748\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__53751\,
            ce => \N__35458\,
            sr => \N__53379\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35602\,
            in1 => \N__34741\,
            in2 => \_gnd_net_\,
            in3 => \N__34724\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__53746\,
            ce => \N__35475\,
            sr => \N__53385\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35618\,
            in1 => \N__34717\,
            in2 => \_gnd_net_\,
            in3 => \N__34700\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__53746\,
            ce => \N__35475\,
            sr => \N__53385\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35599\,
            in1 => \N__34693\,
            in2 => \_gnd_net_\,
            in3 => \N__34676\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__53746\,
            ce => \N__35475\,
            sr => \N__53385\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35615\,
            in1 => \N__35071\,
            in2 => \_gnd_net_\,
            in3 => \N__35054\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__53746\,
            ce => \N__35475\,
            sr => \N__53385\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35600\,
            in1 => \N__35047\,
            in2 => \_gnd_net_\,
            in3 => \N__35030\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__53746\,
            ce => \N__35475\,
            sr => \N__53385\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35616\,
            in1 => \N__35023\,
            in2 => \_gnd_net_\,
            in3 => \N__35006\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__53746\,
            ce => \N__35475\,
            sr => \N__53385\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35601\,
            in1 => \N__34999\,
            in2 => \_gnd_net_\,
            in3 => \N__34982\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__53746\,
            ce => \N__35475\,
            sr => \N__53385\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35617\,
            in1 => \N__34975\,
            in2 => \_gnd_net_\,
            in3 => \N__34958\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__53746\,
            ce => \N__35475\,
            sr => \N__53385\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35603\,
            in1 => \N__34951\,
            in2 => \_gnd_net_\,
            in3 => \N__34934\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_12_21_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__53741\,
            ce => \N__35482\,
            sr => \N__53391\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35611\,
            in1 => \N__34927\,
            in2 => \_gnd_net_\,
            in3 => \N__34910\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__53741\,
            ce => \N__35482\,
            sr => \N__53391\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35604\,
            in1 => \N__34903\,
            in2 => \_gnd_net_\,
            in3 => \N__34886\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__53741\,
            ce => \N__35482\,
            sr => \N__53391\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35612\,
            in1 => \N__35257\,
            in2 => \_gnd_net_\,
            in3 => \N__35240\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__53741\,
            ce => \N__35482\,
            sr => \N__53391\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35605\,
            in1 => \N__35233\,
            in2 => \_gnd_net_\,
            in3 => \N__35216\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__53741\,
            ce => \N__35482\,
            sr => \N__53391\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35613\,
            in1 => \N__35209\,
            in2 => \_gnd_net_\,
            in3 => \N__35192\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__53741\,
            ce => \N__35482\,
            sr => \N__53391\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35606\,
            in1 => \N__35185\,
            in2 => \_gnd_net_\,
            in3 => \N__35168\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__53741\,
            ce => \N__35482\,
            sr => \N__53391\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35614\,
            in1 => \N__35161\,
            in2 => \_gnd_net_\,
            in3 => \N__35144\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__53741\,
            ce => \N__35482\,
            sr => \N__53391\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35607\,
            in1 => \N__35137\,
            in2 => \_gnd_net_\,
            in3 => \N__35120\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_12_22_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__53736\,
            ce => \N__35483\,
            sr => \N__53401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35619\,
            in1 => \N__35113\,
            in2 => \_gnd_net_\,
            in3 => \N__35096\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__53736\,
            ce => \N__35483\,
            sr => \N__53401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35608\,
            in1 => \N__35093\,
            in2 => \_gnd_net_\,
            in3 => \N__35078\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__53736\,
            ce => \N__35483\,
            sr => \N__53401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35620\,
            in1 => \N__35662\,
            in2 => \_gnd_net_\,
            in3 => \N__35645\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__53736\,
            ce => \N__35483\,
            sr => \N__53401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35609\,
            in1 => \N__35641\,
            in2 => \_gnd_net_\,
            in3 => \N__35627\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__53736\,
            ce => \N__35483\,
            sr => \N__53401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__35495\,
            in1 => \N__35610\,
            in2 => \_gnd_net_\,
            in3 => \N__35498\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53736\,
            ce => \N__35483\,
            sr => \N__53401\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35441\,
            in2 => \N__35420\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_16\,
            ltout => OPEN,
            carryin => \bfn_12_23_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15_c_RNIDMOM_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35399\,
            in2 => \N__35381\,
            in3 => \N__35363\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_c_RNIEOPM_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35360\,
            in2 => \N__35342\,
            in3 => \N__35324\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_c_RNIFQQM_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35321\,
            in2 => \N__35303\,
            in3 => \N__35282\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_c_RNIGSRM_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35279\,
            in2 => \N__35981\,
            in3 => \N__35264\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_c_RNIHUSM_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35958\,
            in2 => \N__35849\,
            in3 => \N__35828\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_c_RNI9FMN_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35825\,
            in2 => \N__35982\,
            in3 => \N__35810\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_c_RNIAHNN_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35962\,
            in2 => \N__35807\,
            in3 => \N__35783\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_c_RNIBJON_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35963\,
            in2 => \N__35780\,
            in3 => \N__35762\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_24\,
            ltout => OPEN,
            carryin => \bfn_12_24_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_c_RNICLPN_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35759\,
            in2 => \N__35983\,
            in3 => \N__35741\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_c_RNIDNQN_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35738\,
            in2 => \N__35986\,
            in3 => \N__35723\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_c_RNIEPRN_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35720\,
            in2 => \N__35984\,
            in3 => \N__35705\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_c_RNIFRSN_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35702\,
            in2 => \N__35987\,
            in3 => \N__35687\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_c_RNIGTTN_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35684\,
            in2 => \N__35985\,
            in3 => \N__35669\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_c_RNIHVUN_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35973\,
            in2 => \N__35900\,
            in3 => \N__35882\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35879\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53462\,
            lcout => \GB_BUFFER_red_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35864\,
            in1 => \N__43781\,
            in2 => \_gnd_net_\,
            in3 => \N__40630\,
            lcout => \elapsed_time_ns_1_RNI24CN9_0_15\,
            ltout => \elapsed_time_ns_1_RNI24CN9_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35858\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40631\,
            in1 => \N__44213\,
            in2 => \_gnd_net_\,
            in3 => \N__37729\,
            lcout => \elapsed_time_ns_1_RNI04EN9_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37198\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37351\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35855\,
            in2 => \N__37730\,
            in3 => \N__37483\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36095\,
            in2 => \_gnd_net_\,
            in3 => \N__37471\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37340\,
            in2 => \_gnd_net_\,
            in3 => \N__36089\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38441\,
            in2 => \_gnd_net_\,
            in3 => \N__36074\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36071\,
            in2 => \_gnd_net_\,
            in3 => \N__36053\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37169\,
            in2 => \_gnd_net_\,
            in3 => \N__36038\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37373\,
            in2 => \_gnd_net_\,
            in3 => \N__36023\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37358\,
            in2 => \_gnd_net_\,
            in3 => \N__36008\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37544\,
            in2 => \_gnd_net_\,
            in3 => \N__35990\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37178\,
            in2 => \_gnd_net_\,
            in3 => \N__36227\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37394\,
            in3 => \N__36212\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37421\,
            in2 => \_gnd_net_\,
            in3 => \N__36197\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37490\,
            in2 => \_gnd_net_\,
            in3 => \N__36182\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38366\,
            in2 => \_gnd_net_\,
            in3 => \N__36167\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36164\,
            in2 => \_gnd_net_\,
            in3 => \N__36143\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40493\,
            in2 => \_gnd_net_\,
            in3 => \N__36128\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37565\,
            in2 => \_gnd_net_\,
            in3 => \N__36113\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37559\,
            in2 => \_gnd_net_\,
            in3 => \N__36098\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37415\,
            in2 => \_gnd_net_\,
            in3 => \N__36356\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37427\,
            in2 => \_gnd_net_\,
            in3 => \N__36341\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37508\,
            in2 => \_gnd_net_\,
            in3 => \N__36326\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36323\,
            in2 => \_gnd_net_\,
            in3 => \N__36302\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37529\,
            in2 => \_gnd_net_\,
            in3 => \N__36287\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38492\,
            in2 => \_gnd_net_\,
            in3 => \N__36272\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37553\,
            in2 => \_gnd_net_\,
            in3 => \N__36257\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37451\,
            in3 => \N__36242\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38468\,
            in2 => \_gnd_net_\,
            in3 => \N__36545\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37523\,
            in2 => \_gnd_net_\,
            in3 => \N__36530\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37502\,
            in2 => \_gnd_net_\,
            in3 => \N__36515\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36488\,
            in2 => \_gnd_net_\,
            in3 => \N__36500\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__36497\,
            in1 => \N__37731\,
            in2 => \_gnd_net_\,
            in3 => \N__36491\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38429\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_28_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36478\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53790\,
            ce => \N__37648\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__36467\,
            in1 => \N__36434\,
            in2 => \_gnd_net_\,
            in3 => \N__36397\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__39010\,
            in1 => \N__49750\,
            in2 => \N__39053\,
            in3 => \N__49948\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49946\,
            in1 => \N__38974\,
            in2 => \N__49766\,
            in3 => \N__38990\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__38989\,
            in1 => \N__49944\,
            in2 => \N__38975\,
            in3 => \N__49746\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49945\,
            in1 => \N__39281\,
            in2 => \N__49765\,
            in3 => \N__39301\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__38173\,
            in1 => \N__49751\,
            in2 => \N__38822\,
            in3 => \N__49950\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49947\,
            in1 => \N__38683\,
            in2 => \N__49767\,
            in3 => \N__38037\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__38262\,
            in1 => \N__49752\,
            in2 => \N__38633\,
            in3 => \N__49949\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49951\,
            in1 => \N__38751\,
            in2 => \N__49768\,
            in3 => \N__38317\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49942\,
            in1 => \N__39349\,
            in2 => \N__49757\,
            in3 => \N__38193\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__39350\,
            in1 => \N__49941\,
            in2 => \N__38195\,
            in3 => \N__49712\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39103\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53785\,
            ce => \N__39076\,
            sr => \N__53342\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__38936\,
            in1 => \N__49713\,
            in2 => \N__38906\,
            in3 => \N__49940\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37821\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__36590\,
            in1 => \_gnd_net_\,
            in2 => \N__36566\,
            in3 => \N__49936\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \N__49714\,
            in1 => \N__38902\,
            in2 => \N__50021\,
            in3 => \N__38935\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__36589\,
            in1 => \N__49935\,
            in2 => \_gnd_net_\,
            in3 => \N__36563\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38125\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36582\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__49996\,
            in1 => \N__49553\,
            in2 => \N__38000\,
            in3 => \N__40735\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49554\,
            in1 => \N__49997\,
            in2 => \N__40739\,
            in3 => \N__37999\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__49998\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49552\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39578\,
            in1 => \N__40734\,
            in2 => \_gnd_net_\,
            in3 => \N__37995\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__39577\,
            in1 => \N__37822\,
            in2 => \_gnd_net_\,
            in3 => \N__36583\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39107\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53780\,
            ce => \N__39075\,
            sr => \N__53354\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45227\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53780\,
            ce => \N__39075\,
            sr => \N__53354\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49992\,
            in1 => \N__49717\,
            in2 => \N__38821\,
            in3 => \N__38174\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49719\,
            in1 => \N__49994\,
            in2 => \N__40804\,
            in3 => \N__38214\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38859\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__49715\,
            in1 => \N__49995\,
            in2 => \N__39539\,
            in3 => \N__41273\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39419\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49718\,
            in1 => \N__49993\,
            in2 => \N__39725\,
            in3 => \N__39682\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49991\,
            in1 => \N__49716\,
            in2 => \N__38684\,
            in3 => \N__38039\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__49979\,
            in1 => \N__38146\,
            in2 => \N__45944\,
            in3 => \N__38124\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45191\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53770\,
            ce => \N__39074\,
            sr => \N__53365\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__38147\,
            in1 => \N__49978\,
            in2 => \N__38126\,
            in3 => \N__45943\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__49980\,
            in1 => \N__49623\,
            in2 => \N__46427\,
            in3 => \N__38334\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110011"
        )
    port map (
            in0 => \N__49622\,
            in1 => \N__49981\,
            in2 => \N__38341\,
            in3 => \N__46421\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__39902\,
            in1 => \N__49727\,
            in2 => \N__39389\,
            in3 => \N__49986\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101111"
        )
    port map (
            in0 => \N__39458\,
            in1 => \N__49728\,
            in2 => \N__50141\,
            in3 => \N__39431\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49990\,
            in1 => \N__38866\,
            in2 => \N__49761\,
            in3 => \N__38242\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__38867\,
            in1 => \N__49736\,
            in2 => \N__38243\,
            in3 => \N__49989\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49988\,
            in1 => \N__40805\,
            in2 => \N__49760\,
            in3 => \N__38219\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__38318\,
            in1 => \N__49729\,
            in2 => \N__38759\,
            in3 => \N__49987\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49985\,
            in1 => \N__38625\,
            in2 => \N__49759\,
            in3 => \N__38270\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38533\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38287\,
            ce => 'H',
            sr => \N__53380\
        );

    \pwm_generator_inst.un3_threshold_axb_8_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36812\,
            in2 => \N__36791\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_21_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36758\,
            in2 => \N__36740\,
            in3 => \N__36707\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36704\,
            in2 => \N__36683\,
            in3 => \N__36650\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36647\,
            in2 => \N__36629\,
            in3 => \N__36593\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37163\,
            in2 => \N__36884\,
            in3 => \N__37130\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36866\,
            in2 => \N__37127\,
            in3 => \N__37094\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37091\,
            in2 => \N__36885\,
            in3 => \N__37064\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36870\,
            in2 => \N__37061\,
            in3 => \N__37025\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36886\,
            in2 => \N__37022\,
            in3 => \N__36989\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_13_22_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36986\,
            in2 => \N__36897\,
            in3 => \N__36956\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36953\,
            in2 => \N__36899\,
            in3 => \N__36920\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36917\,
            in2 => \N__36898\,
            in3 => \N__37322\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_LUT4_0_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37319\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__53461\,
            in1 => \N__37300\,
            in2 => \_gnd_net_\,
            in3 => \N__37231\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37304\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53738\,
            ce => 'H',
            sr => \N__53402\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40225\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53738\,
            ce => 'H',
            sr => \N__53402\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__40156\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53738\,
            ce => 'H',
            sr => \N__53402\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40605\,
            in1 => \N__37199\,
            in2 => \_gnd_net_\,
            in3 => \N__44000\,
            lcout => \elapsed_time_ns_1_RNI03DN9_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37187\,
            in1 => \N__43889\,
            in2 => \_gnd_net_\,
            in3 => \N__40604\,
            lcout => \elapsed_time_ns_1_RNITUBN9_0_10\,
            ltout => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37181\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38386\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37403\,
            in1 => \N__43865\,
            in2 => \_gnd_net_\,
            in3 => \N__40582\,
            lcout => \elapsed_time_ns_1_RNIUVBN9_0_11\,
            ltout => \elapsed_time_ns_1_RNIUVBN9_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37397\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43612\,
            in1 => \N__37382\,
            in2 => \_gnd_net_\,
            in3 => \N__40580\,
            lcout => \elapsed_time_ns_1_RNIJ53T9_0_7\,
            ltout => \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37376\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37367\,
            in1 => \N__43583\,
            in2 => \_gnd_net_\,
            in3 => \N__40581\,
            lcout => \elapsed_time_ns_1_RNIK63T9_0_8\,
            ltout => \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37361\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37352\,
            in1 => \N__40583\,
            in2 => \_gnd_net_\,
            in3 => \N__43655\,
            lcout => \elapsed_time_ns_1_RNIH33T9_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38398\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38581\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37484\,
            in1 => \N__40409\,
            in2 => \_gnd_net_\,
            in3 => \N__40619\,
            lcout => \elapsed_time_ns_1_RNIDV2T9_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40620\,
            in1 => \N__37472\,
            in2 => \_gnd_net_\,
            in3 => \N__40391\,
            lcout => \elapsed_time_ns_1_RNIE03T9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37439\,
            in1 => \N__44042\,
            in2 => \_gnd_net_\,
            in3 => \N__40621\,
            lcout => \elapsed_time_ns_1_RNIU0DN9_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37460\,
            in1 => \N__43910\,
            in2 => \_gnd_net_\,
            in3 => \N__40618\,
            lcout => \elapsed_time_ns_1_RNI47DN9_0_26\,
            ltout => \elapsed_time_ns_1_RNI47DN9_0_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37454\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37438\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38353\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40622\,
            in1 => \N__37409\,
            in2 => \_gnd_net_\,
            in3 => \N__43556\,
            lcout => \elapsed_time_ns_1_RNIL73T9_0_9\,
            ltout => \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37547\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37538\,
            in1 => \N__43979\,
            in2 => \_gnd_net_\,
            in3 => \N__40623\,
            lcout => \elapsed_time_ns_1_RNI14DN9_0_23\,
            ltout => \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37532\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38455\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40625\,
            in1 => \N__37517\,
            in2 => \_gnd_net_\,
            in3 => \N__44021\,
            lcout => \elapsed_time_ns_1_RNIV1DN9_0_21\,
            ltout => \elapsed_time_ns_1_RNIV1DN9_0_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37511\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40649\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37496\,
            in1 => \N__43742\,
            in2 => \_gnd_net_\,
            in3 => \N__40624\,
            lcout => \elapsed_time_ns_1_RNI46CN9_0_17\,
            ltout => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37568\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38512\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38704\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38604\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38952\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38655\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39032\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38730\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41696\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39263\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42828\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__50059\,
            in1 => \N__40851\,
            in2 => \N__49769\,
            in3 => \N__38092\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49785\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39738\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38922\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_0_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37736\,
            in2 => \_gnd_net_\,
            in3 => \N__37685\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53791\,
            ce => \N__37643\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41801\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38790\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39190\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39363\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39495\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39699\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39129\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37829\,
            in2 => \N__37823\,
            in3 => \N__37820\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37796\,
            in2 => \_gnd_net_\,
            in3 => \N__37787\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37784\,
            in2 => \_gnd_net_\,
            in3 => \N__37775\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37772\,
            in2 => \_gnd_net_\,
            in3 => \N__37763\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37760\,
            in2 => \_gnd_net_\,
            in3 => \N__37751\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37748\,
            in2 => \_gnd_net_\,
            in3 => \N__37739\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37919\,
            in2 => \_gnd_net_\,
            in3 => \N__37910\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37907\,
            in2 => \_gnd_net_\,
            in3 => \N__37898\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39317\,
            in2 => \_gnd_net_\,
            in3 => \N__37895\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37892\,
            in2 => \_gnd_net_\,
            in3 => \N__37883\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37880\,
            in2 => \_gnd_net_\,
            in3 => \N__37871\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37868\,
            in2 => \_gnd_net_\,
            in3 => \N__37859\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37856\,
            in2 => \_gnd_net_\,
            in3 => \N__37844\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37841\,
            in2 => \_gnd_net_\,
            in3 => \N__37832\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40829\,
            in2 => \_gnd_net_\,
            in3 => \N__38018\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38015\,
            in2 => \_gnd_net_\,
            in3 => \N__38006\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40751\,
            in2 => \_gnd_net_\,
            in3 => \N__38003\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40709\,
            in2 => \_gnd_net_\,
            in3 => \N__37985\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37982\,
            in2 => \_gnd_net_\,
            in3 => \N__37970\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37967\,
            in2 => \_gnd_net_\,
            in3 => \N__37958\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37955\,
            in2 => \_gnd_net_\,
            in3 => \N__37946\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37943\,
            in2 => \_gnd_net_\,
            in3 => \N__37934\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37931\,
            in2 => \_gnd_net_\,
            in3 => \N__37922\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40817\,
            in2 => \_gnd_net_\,
            in3 => \N__38072\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40763\,
            in2 => \_gnd_net_\,
            in3 => \N__38069\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38066\,
            in2 => \_gnd_net_\,
            in3 => \N__38060\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40697\,
            in2 => \_gnd_net_\,
            in3 => \N__38057\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41237\,
            in2 => \_gnd_net_\,
            in3 => \N__38054\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38051\,
            in2 => \_gnd_net_\,
            in3 => \N__38045\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38042\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__49639\,
            in1 => \N__50049\,
            in2 => \N__38096\,
            in3 => \N__40861\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39585\,
            in1 => \N__38673\,
            in2 => \_gnd_net_\,
            in3 => \N__38038\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__39481\,
            in1 => \N__50096\,
            in2 => \N__49758\,
            in3 => \N__39515\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__50095\,
            in1 => \N__49723\,
            in2 => \N__39218\,
            in3 => \N__39241\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39348\,
            in1 => \N__39653\,
            in2 => \_gnd_net_\,
            in3 => \N__38194\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__39657\,
            in1 => \_gnd_net_\,
            in2 => \N__41722\,
            in3 => \N__41745\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__38808\,
            in1 => \N__39655\,
            in2 => \_gnd_net_\,
            in3 => \N__38172\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39656\,
            in1 => \N__39754\,
            in2 => \_gnd_net_\,
            in3 => \N__39778\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__38140\,
            in1 => \N__38120\,
            in2 => \_gnd_net_\,
            in3 => \N__39652\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__39654\,
            in1 => \_gnd_net_\,
            in2 => \N__42850\,
            in3 => \N__42876\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__39635\,
            in1 => \_gnd_net_\,
            in2 => \N__40862\,
            in3 => \N__38091\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39214\,
            in1 => \N__39637\,
            in2 => \_gnd_net_\,
            in3 => \N__39240\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39633\,
            in1 => \N__38629\,
            in2 => \_gnd_net_\,
            in3 => \N__38269\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41820\,
            in1 => \N__39636\,
            in2 => \_gnd_net_\,
            in3 => \N__41776\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__39639\,
            in1 => \N__39174\,
            in2 => \_gnd_net_\,
            in3 => \N__39147\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39381\,
            in1 => \N__39634\,
            in2 => \_gnd_net_\,
            in3 => \N__39901\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39638\,
            in1 => \N__39513\,
            in2 => \_gnd_net_\,
            in3 => \N__39480\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__50118\,
            in1 => \N__38865\,
            in2 => \_gnd_net_\,
            in3 => \N__38238\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42987\,
            in1 => \N__39664\,
            in2 => \_gnd_net_\,
            in3 => \N__42943\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__50117\,
            in1 => \N__40797\,
            in2 => \_gnd_net_\,
            in3 => \N__38215\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39430\,
            in1 => \N__50121\,
            in2 => \_gnd_net_\,
            in3 => \N__39451\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111000101"
        )
    port map (
            in0 => \N__39148\,
            in1 => \N__39179\,
            in2 => \N__50135\,
            in3 => \N__49624\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41272\,
            in1 => \N__50120\,
            in2 => \_gnd_net_\,
            in3 => \N__39538\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__41674\,
            in1 => \_gnd_net_\,
            in2 => \N__39665\,
            in3 => \N__41634\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50119\,
            in2 => \N__43066\,
            in3 => \N__43107\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50091\,
            in2 => \_gnd_net_\,
            in3 => \N__38342\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__38310\,
            in1 => \N__39660\,
            in2 => \_gnd_net_\,
            in3 => \N__38752\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38532\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38288\,
            ce => 'H',
            sr => \N__53381\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__43582\,
            in1 => \N__40421\,
            in2 => \N__43613\,
            in3 => \N__40415\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43676\,
            in1 => \N__38276\,
            in2 => \_gnd_net_\,
            in3 => \N__40577\,
            lcout => \elapsed_time_ns_1_RNIG23T9_0_4\,
            ltout => \elapsed_time_ns_1_RNIG23T9_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38444\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44234\,
            in1 => \N__38425\,
            in2 => \_gnd_net_\,
            in3 => \N__40579\,
            lcout => \elapsed_time_ns_1_RNIV2EN9_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40679\,
            in1 => \N__40664\,
            in2 => \N__40658\,
            in3 => \N__40685\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__44209\,
            in1 => \N__40670\,
            in2 => \N__38411\,
            in3 => \N__38408\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__38399\,
            in1 => \_gnd_net_\,
            in2 => \N__38402\,
            in3 => \N__43694\,
            lcout => \elapsed_time_ns_1_RNIF13T9_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38387\,
            in1 => \N__43634\,
            in2 => \_gnd_net_\,
            in3 => \N__40578\,
            lcout => \elapsed_time_ns_1_RNII43T9_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43802\,
            in1 => \N__38375\,
            in2 => \_gnd_net_\,
            in3 => \N__40606\,
            lcout => \elapsed_time_ns_1_RNI13CN9_0_14\,
            ltout => \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38369\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40607\,
            in1 => \N__38354\,
            in2 => \_gnd_net_\,
            in3 => \N__43844\,
            lcout => \elapsed_time_ns_1_RNIV0CN9_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40610\,
            in1 => \N__38480\,
            in2 => \_gnd_net_\,
            in3 => \N__44291\,
            lcout => \elapsed_time_ns_1_RNI58DN9_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38582\,
            in1 => \N__43823\,
            in2 => \_gnd_net_\,
            in3 => \N__40608\,
            lcout => \elapsed_time_ns_1_RNI02CN9_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40609\,
            in1 => \N__38570\,
            in2 => \_gnd_net_\,
            in3 => \N__44063\,
            lcout => \elapsed_time_ns_1_RNI68CN9_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__41105\,
            in1 => \N__38551\,
            in2 => \_gnd_net_\,
            in3 => \N__41141\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_166_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40627\,
            in1 => \N__38513\,
            in2 => \_gnd_net_\,
            in3 => \N__43718\,
            lcout => \elapsed_time_ns_1_RNI57CN9_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38501\,
            in1 => \N__43955\,
            in2 => \_gnd_net_\,
            in3 => \N__40626\,
            lcout => \elapsed_time_ns_1_RNI25DN9_0_24\,
            ltout => \elapsed_time_ns_1_RNI25DN9_0_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38495\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38479\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40629\,
            in1 => \N__38456\,
            in2 => \_gnd_net_\,
            in3 => \N__44270\,
            lcout => \elapsed_time_ns_1_RNI69DN9_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38705\,
            in1 => \N__43934\,
            in2 => \_gnd_net_\,
            in3 => \N__40628\,
            lcout => \elapsed_time_ns_1_RNI36DN9_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45151\,
            in2 => \N__45223\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__53814\,
            ce => \N__39080\,
            sr => \N__53327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45127\,
            in2 => \N__45190\,
            in3 => \N__38693\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__53814\,
            ce => \N__39080\,
            sr => \N__53327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45152\,
            in2 => \N__45103\,
            in3 => \N__38690\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__53814\,
            ce => \N__39080\,
            sr => \N__53327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45128\,
            in2 => \N__45073\,
            in3 => \N__38687\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__53814\,
            ce => \N__39080\,
            sr => \N__53327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45040\,
            in2 => \N__45104\,
            in3 => \N__38639\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__53814\,
            ce => \N__39080\,
            sr => \N__53327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45643\,
            in2 => \N__45074\,
            in3 => \N__38636\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__53814\,
            ce => \N__39080\,
            sr => \N__53327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45616\,
            in2 => \N__45044\,
            in3 => \N__38588\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__53814\,
            ce => \N__39080\,
            sr => \N__53327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45644\,
            in2 => \N__45583\,
            in3 => \N__38585\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__53814\,
            ce => \N__39080\,
            sr => \N__53327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45541\,
            in2 => \N__45620\,
            in3 => \N__38825\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__53805\,
            ce => \N__39079\,
            sr => \N__53329\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45514\,
            in2 => \N__45584\,
            in3 => \N__38774\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__53805\,
            ce => \N__39079\,
            sr => \N__53329\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45490\,
            in2 => \N__45545\,
            in3 => \N__38771\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__53805\,
            ce => \N__39079\,
            sr => \N__53329\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45515\,
            in2 => \N__45466\,
            in3 => \N__38768\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__53805\,
            ce => \N__39079\,
            sr => \N__53329\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45491\,
            in2 => \N__45436\,
            in3 => \N__38765\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__53805\,
            ce => \N__39079\,
            sr => \N__53329\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45910\,
            in2 => \N__45467\,
            in3 => \N__38762\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__53805\,
            ce => \N__39079\,
            sr => \N__53329\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45883\,
            in2 => \N__45437\,
            in3 => \N__38714\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__53805\,
            ce => \N__39079\,
            sr => \N__53329\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45911\,
            in2 => \N__45850\,
            in3 => \N__38711\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__53805\,
            ce => \N__39079\,
            sr => \N__53329\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45808\,
            in2 => \N__45887\,
            in3 => \N__38708\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__53799\,
            ce => \N__39078\,
            sr => \N__53335\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45781\,
            in2 => \N__45851\,
            in3 => \N__38888\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__53799\,
            ce => \N__39078\,
            sr => \N__53335\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45754\,
            in2 => \N__45812\,
            in3 => \N__38885\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__53799\,
            ce => \N__39078\,
            sr => \N__53335\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45782\,
            in2 => \N__45727\,
            in3 => \N__38882\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__53799\,
            ce => \N__39078\,
            sr => \N__53335\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45694\,
            in2 => \N__45758\,
            in3 => \N__38879\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__53799\,
            ce => \N__39078\,
            sr => \N__53335\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45667\,
            in2 => \N__45728\,
            in3 => \N__38876\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__53799\,
            ce => \N__39078\,
            sr => \N__53335\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46165\,
            in2 => \N__45698\,
            in3 => \N__38873\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__53799\,
            ce => \N__39078\,
            sr => \N__53335\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45668\,
            in2 => \N__46132\,
            in3 => \N__38870\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__53799\,
            ce => \N__39078\,
            sr => \N__53335\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46093\,
            in2 => \N__46169\,
            in3 => \N__38831\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__53792\,
            ce => \N__39077\,
            sr => \N__53337\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46069\,
            in2 => \N__46133\,
            in3 => \N__38828\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__53792\,
            ce => \N__39077\,
            sr => \N__53337\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46094\,
            in2 => \N__46046\,
            in3 => \N__39116\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__53792\,
            ce => \N__39077\,
            sr => \N__53337\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46070\,
            in2 => \N__46016\,
            in3 => \N__39113\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__53792\,
            ce => \N__39077\,
            sr => \N__53337\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39110\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39096\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53792\,
            ce => \N__39077\,
            sr => \N__53337\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39280\,
            in1 => \N__39649\,
            in2 => \_gnd_net_\,
            in3 => \N__39297\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39651\,
            in1 => \N__39042\,
            in2 => \_gnd_net_\,
            in3 => \N__39006\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__38988\,
            in1 => \N__39650\,
            in2 => \_gnd_net_\,
            in3 => \N__38965\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39648\,
            in1 => \N__38929\,
            in2 => \_gnd_net_\,
            in3 => \N__38901\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \N__49649\,
            in1 => \N__39777\,
            in2 => \N__50126\,
            in3 => \N__39753\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__41749\,
            in1 => \N__50111\,
            in2 => \N__41723\,
            in3 => \N__49650\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39339\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39311\,
            in1 => \_gnd_net_\,
            in2 => \N__42703\,
            in3 => \N__39872\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49558\,
            in1 => \N__50089\,
            in2 => \N__39724\,
            in3 => \N__39683\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__50087\,
            in1 => \N__49559\,
            in2 => \N__41821\,
            in3 => \N__41775\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__49555\,
            in1 => \N__50083\,
            in2 => \N__39305\,
            in3 => \N__39279\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__50086\,
            in1 => \N__41670\,
            in2 => \N__41638\,
            in3 => \N__49563\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__49561\,
            in1 => \N__50088\,
            in2 => \N__39242\,
            in3 => \N__39213\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__50090\,
            in1 => \N__49560\,
            in2 => \N__39178\,
            in3 => \N__39149\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__49557\,
            in1 => \N__50085\,
            in2 => \N__39779\,
            in3 => \N__39755\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__50084\,
            in1 => \N__49556\,
            in2 => \N__42880\,
            in3 => \N__42843\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39658\,
            in1 => \N__49792\,
            in2 => \_gnd_net_\,
            in3 => \N__50158\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__39708\,
            in1 => \N__39681\,
            in2 => \_gnd_net_\,
            in3 => \N__39659\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42991\,
            in1 => \N__50099\,
            in2 => \N__49708\,
            in3 => \N__42942\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__50101\,
            in1 => \N__41268\,
            in2 => \N__49706\,
            in3 => \N__39537\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__39514\,
            in1 => \N__50098\,
            in2 => \N__39482\,
            in3 => \N__49634\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__50100\,
            in1 => \N__43108\,
            in2 => \N__49705\,
            in3 => \N__43059\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__39450\,
            in1 => \N__49635\,
            in2 => \N__39429\,
            in3 => \N__50102\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__50097\,
            in1 => \N__39385\,
            in2 => \N__49707\,
            in3 => \N__39897\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39871\,
            in2 => \N__46419\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42416\,
            in2 => \N__39848\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39836\,
            in2 => \N__42549\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42420\,
            in2 => \N__39827\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39818\,
            in2 => \N__42550\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42424\,
            in2 => \N__39809\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39797\,
            in2 => \N__42551\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42428\,
            in2 => \N__39791\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42542\,
            in2 => \N__39962\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39953\,
            in2 => \N__42623\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42530\,
            in2 => \N__39947\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39938\,
            in2 => \N__42620\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42534\,
            in2 => \N__39932\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39923\,
            in2 => \N__42621\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42538\,
            in2 => \N__39917\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39908\,
            in2 => \N__42622\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42514\,
            in2 => \N__40049\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40037\,
            in2 => \N__42616\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42518\,
            in2 => \N__40031\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40013\,
            in2 => \N__42617\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42522\,
            in2 => \N__40007\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39998\,
            in2 => \N__42618\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42526\,
            in2 => \N__39992\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39977\,
            in2 => \N__42619\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42501\,
            in2 => \N__39971\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40103\,
            in2 => \N__42613\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42505\,
            in2 => \N__40097\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40088\,
            in2 => \N__42614\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42509\,
            in2 => \N__40082\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40073\,
            in2 => \N__42615\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42513\,
            in2 => \N__40067\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50125\,
            in2 => \_gnd_net_\,
            in3 => \N__40058\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40055\,
            in2 => \_gnd_net_\,
            in3 => \N__46805\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47159\,
            in2 => \_gnd_net_\,
            in3 => \N__40130\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__53759\,
            ce => 'H',
            sr => \N__53374\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47138\,
            in2 => \_gnd_net_\,
            in3 => \N__40127\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__53759\,
            ce => 'H',
            sr => \N__53374\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47117\,
            in2 => \_gnd_net_\,
            in3 => \N__40124\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__53759\,
            ce => 'H',
            sr => \N__53374\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47096\,
            in2 => \_gnd_net_\,
            in3 => \N__40121\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__53759\,
            ce => 'H',
            sr => \N__53374\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47075\,
            in2 => \_gnd_net_\,
            in3 => \N__40118\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__53759\,
            ce => 'H',
            sr => \N__53374\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47054\,
            in2 => \_gnd_net_\,
            in3 => \N__40115\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__53759\,
            ce => 'H',
            sr => \N__53374\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47033\,
            in2 => \_gnd_net_\,
            in3 => \N__40112\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__53759\,
            ce => 'H',
            sr => \N__53374\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47012\,
            in2 => \_gnd_net_\,
            in3 => \N__40109\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__53753\,
            ce => 'H',
            sr => \N__53382\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47339\,
            in2 => \_gnd_net_\,
            in3 => \N__40106\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__53753\,
            ce => 'H',
            sr => \N__53382\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47318\,
            in2 => \_gnd_net_\,
            in3 => \N__40181\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__53753\,
            ce => 'H',
            sr => \N__53382\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47297\,
            in2 => \_gnd_net_\,
            in3 => \N__40178\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__53753\,
            ce => 'H',
            sr => \N__53382\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47273\,
            in2 => \_gnd_net_\,
            in3 => \N__40175\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__53753\,
            ce => 'H',
            sr => \N__53382\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47249\,
            in2 => \_gnd_net_\,
            in3 => \N__40172\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__53753\,
            ce => 'H',
            sr => \N__53382\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47225\,
            in2 => \_gnd_net_\,
            in3 => \N__40169\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            clk => \N__53753\,
            ce => 'H',
            sr => \N__53382\
        );

    \current_shift_inst.PI_CTRL.error_control_15_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47204\,
            in2 => \_gnd_net_\,
            in3 => \N__40166\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            clk => \N__53753\,
            ce => 'H',
            sr => \N__53382\
        );

    \current_shift_inst.PI_CTRL.error_control_16_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47180\,
            in2 => \_gnd_net_\,
            in3 => \N__40163\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_16\,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            clk => \N__53748\,
            ce => 'H',
            sr => \N__53386\
        );

    \current_shift_inst.PI_CTRL.error_control_17_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47513\,
            in2 => \_gnd_net_\,
            in3 => \N__40136\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            clk => \N__53748\,
            ce => 'H',
            sr => \N__53386\
        );

    \current_shift_inst.PI_CTRL.error_control_18_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47486\,
            in2 => \_gnd_net_\,
            in3 => \N__40133\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            clk => \N__53748\,
            ce => 'H',
            sr => \N__53386\
        );

    \current_shift_inst.PI_CTRL.error_control_19_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47459\,
            in2 => \_gnd_net_\,
            in3 => \N__40208\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            clk => \N__53748\,
            ce => 'H',
            sr => \N__53386\
        );

    \current_shift_inst.PI_CTRL.error_control_20_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47438\,
            in2 => \_gnd_net_\,
            in3 => \N__40205\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            clk => \N__53748\,
            ce => 'H',
            sr => \N__53386\
        );

    \current_shift_inst.PI_CTRL.error_control_21_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47417\,
            in2 => \_gnd_net_\,
            in3 => \N__40202\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            clk => \N__53748\,
            ce => 'H',
            sr => \N__53386\
        );

    \current_shift_inst.PI_CTRL.error_control_22_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47393\,
            in2 => \_gnd_net_\,
            in3 => \N__40199\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            clk => \N__53748\,
            ce => 'H',
            sr => \N__53386\
        );

    \current_shift_inst.PI_CTRL.error_control_23_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47372\,
            in2 => \_gnd_net_\,
            in3 => \N__40196\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            clk => \N__53748\,
            ce => 'H',
            sr => \N__53386\
        );

    \current_shift_inst.PI_CTRL.error_control_24_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47831\,
            in2 => \_gnd_net_\,
            in3 => \N__40193\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_24\,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            clk => \N__53743\,
            ce => 'H',
            sr => \N__53392\
        );

    \current_shift_inst.PI_CTRL.error_control_25_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47810\,
            in2 => \_gnd_net_\,
            in3 => \N__40190\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            clk => \N__53743\,
            ce => 'H',
            sr => \N__53392\
        );

    \current_shift_inst.PI_CTRL.error_control_26_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47783\,
            in2 => \_gnd_net_\,
            in3 => \N__40187\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            clk => \N__53743\,
            ce => 'H',
            sr => \N__53392\
        );

    \current_shift_inst.PI_CTRL.error_control_27_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47762\,
            in2 => \_gnd_net_\,
            in3 => \N__40184\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            clk => \N__53743\,
            ce => 'H',
            sr => \N__53392\
        );

    \current_shift_inst.PI_CTRL.error_control_28_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47738\,
            in2 => \_gnd_net_\,
            in3 => \N__40370\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            clk => \N__53743\,
            ce => 'H',
            sr => \N__53392\
        );

    \current_shift_inst.PI_CTRL.error_control_29_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47723\,
            in2 => \_gnd_net_\,
            in3 => \N__40367\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            clk => \N__53743\,
            ce => 'H',
            sr => \N__53392\
        );

    \current_shift_inst.PI_CTRL.error_control_30_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43397\,
            in2 => \_gnd_net_\,
            in3 => \N__40364\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_30\,
            clk => \N__53743\,
            ce => 'H',
            sr => \N__53392\
        );

    \current_shift_inst.PI_CTRL.error_control_31_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47705\,
            in2 => \_gnd_net_\,
            in3 => \N__40361\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53743\,
            ce => 'H',
            sr => \N__53392\
        );

    \current_shift_inst.PI_CTRL.prop_term_30_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40351\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53739\,
            ce => 'H',
            sr => \N__53403\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40327\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53739\,
            ce => 'H',
            sr => \N__53403\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40300\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53739\,
            ce => 'H',
            sr => \N__53403\
        );

    \current_shift_inst.PI_CTRL.prop_term_29_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40273\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53739\,
            ce => 'H',
            sr => \N__53403\
        );

    \current_shift_inst.PI_CTRL.prop_term_27_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40255\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53732\,
            ce => 'H',
            sr => \N__53407\
        );

    \current_shift_inst.PI_CTRL.prop_term_26_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40474\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53732\,
            ce => 'H',
            sr => \N__53407\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40450\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53732\,
            ce => 'H',
            sr => \N__53407\
        );

    \current_shift_inst.PI_CTRL.prop_term_31_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40430\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53732\,
            ce => 'H',
            sr => \N__53407\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52423\,
            in1 => \N__48188\,
            in2 => \_gnd_net_\,
            in3 => \N__52240\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53730\,
            ce => 'H',
            sr => \N__53411\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_15_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__52417\,
            in1 => \N__52196\,
            in2 => \_gnd_net_\,
            in3 => \N__48350\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53728\,
            ce => 'H',
            sr => \N__53414\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_15_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52416\,
            in1 => \N__48134\,
            in2 => \_gnd_net_\,
            in3 => \N__52197\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53728\,
            ce => 'H',
            sr => \N__53414\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43687\,
            in1 => \N__43669\,
            in2 => \N__40387\,
            in3 => \N__40402\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__43627\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43648\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_16_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__44150\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53852\,
            ce => \N__44192\,
            sr => \N__53314\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_16_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__44119\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53852\,
            ce => \N__44192\,
            sr => \N__53314\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43774\,
            in1 => \N__43732\,
            in2 => \N__43714\,
            in3 => \N__43756\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44014\,
            in1 => \N__44035\,
            in2 => \N__43999\,
            in3 => \N__44056\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43885\,
            in1 => \N__43858\,
            in2 => \N__43552\,
            in3 => \N__43837\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43795\,
            in2 => \N__40673\,
            in3 => \N__43816\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44248\,
            in1 => \N__43948\,
            in2 => \N__43975\,
            in3 => \N__44230\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44284\,
            in1 => \N__43903\,
            in2 => \N__43930\,
            in3 => \N__44263\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40617\,
            in1 => \N__40645\,
            in2 => \_gnd_net_\,
            in3 => \N__44249\,
            lcout => \elapsed_time_ns_1_RNI7ADN9_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40502\,
            in1 => \N__43760\,
            in2 => \_gnd_net_\,
            in3 => \N__40616\,
            lcout => \elapsed_time_ns_1_RNI35CN9_0_16\,
            ltout => \elapsed_time_ns_1_RNI35CN9_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40496\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41104\,
            in2 => \_gnd_net_\,
            in3 => \N__41140\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_165_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41103\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_0_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41078\,
            in2 => \_gnd_net_\,
            in3 => \N__41021\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53806\,
            ce => \N__40967\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40845\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42968\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40779\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41657\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40720\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43088\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41255\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42796\,
            in2 => \N__45983\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_13_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45931\,
            in2 => \N__41225\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49487\,
            in2 => \N__41207\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49157\,
            in2 => \N__49612\,
            in3 => \N__41195\,
            lcout => \current_shift_inst.un38_control_input_0_s1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49491\,
            in2 => \N__41192\,
            in3 => \N__41180\,
            lcout => \current_shift_inst.un38_control_input_0_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41177\,
            in2 => \N__49613\,
            in3 => \N__41165\,
            lcout => \current_shift_inst.un38_control_input_0_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49495\,
            in2 => \N__41162\,
            in3 => \N__41144\,
            lcout => \current_shift_inst.un38_control_input_0_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41393\,
            in2 => \N__49614\,
            in3 => \N__41384\,
            lcout => \current_shift_inst.un38_control_input_0_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49326\,
            in2 => \N__41381\,
            in3 => \N__41363\,
            lcout => \current_shift_inst.un38_control_input_0_s1_8\,
            ltout => OPEN,
            carryin => \bfn_16_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41360\,
            in2 => \N__49502\,
            in3 => \N__41348\,
            lcout => \current_shift_inst.un38_control_input_0_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49330\,
            in2 => \N__42812\,
            in3 => \N__41345\,
            lcout => \current_shift_inst.un38_control_input_0_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41342\,
            in2 => \N__49503\,
            in3 => \N__41330\,
            lcout => \current_shift_inst.un38_control_input_0_s1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49334\,
            in2 => \N__41327\,
            in3 => \N__41312\,
            lcout => \current_shift_inst.un38_control_input_0_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41309\,
            in2 => \N__49504\,
            in3 => \N__41303\,
            lcout => \current_shift_inst.un38_control_input_0_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49338\,
            in2 => \N__41300\,
            in3 => \N__41291\,
            lcout => \current_shift_inst.un38_control_input_0_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41288\,
            in2 => \N__49505\,
            in3 => \N__41276\,
            lcout => \current_shift_inst.un38_control_input_0_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49404\,
            in2 => \N__41486\,
            in3 => \N__41471\,
            lcout => \current_shift_inst.un38_control_input_0_s1_16\,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41468\,
            in2 => \N__49545\,
            in3 => \N__41462\,
            lcout => \current_shift_inst.un38_control_input_0_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49408\,
            in2 => \N__41459\,
            in3 => \N__41447\,
            lcout => \current_shift_inst.un38_control_input_0_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41444\,
            in2 => \N__49546\,
            in3 => \N__41438\,
            lcout => \current_shift_inst.un38_control_input_0_s1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49412\,
            in2 => \N__41435\,
            in3 => \N__41426\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41423\,
            in2 => \N__49547\,
            in3 => \N__41417\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49416\,
            in2 => \N__41414\,
            in3 => \N__41405\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41402\,
            in2 => \N__49548\,
            in3 => \N__41396\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49420\,
            in2 => \N__41591\,
            in3 => \N__41582\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41579\,
            in2 => \N__49549\,
            in3 => \N__41567\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49424\,
            in2 => \N__41564\,
            in3 => \N__41549\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41546\,
            in2 => \N__49550\,
            in3 => \N__41540\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49428\,
            in2 => \N__41537\,
            in3 => \N__41528\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41525\,
            in2 => \N__49551\,
            in3 => \N__41519\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49432\,
            in2 => \N__41516\,
            in3 => \N__41501\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__49433\,
            in1 => \N__50103\,
            in2 => \_gnd_net_\,
            in3 => \N__41498\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__41495\,
            in1 => \N__46706\,
            in2 => \_gnd_net_\,
            in3 => \N__47680\,
            lcout => \current_shift_inst.control_input_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__50104\,
            in1 => \N__49539\,
            in2 => \N__42887\,
            in3 => \N__42851\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__42800\,
            in1 => \N__42552\,
            in2 => \_gnd_net_\,
            in3 => \N__46420\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__41831\,
            in1 => \N__46898\,
            in2 => \_gnd_net_\,
            in3 => \N__47681\,
            lcout => \current_shift_inst.control_input_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__50107\,
            in1 => \N__49540\,
            in2 => \N__41825\,
            in3 => \N__41780\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__49541\,
            in1 => \N__50105\,
            in2 => \N__41753\,
            in3 => \N__41718\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__50106\,
            in1 => \N__49542\,
            in2 => \N__41678\,
            in3 => \N__41639\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__47663\,
            in1 => \N__41609\,
            in2 => \_gnd_net_\,
            in3 => \N__46943\,
            lcout => \current_shift_inst.control_input_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__47671\,
            in1 => \N__41600\,
            in2 => \_gnd_net_\,
            in3 => \N__46682\,
            lcout => \current_shift_inst.control_input_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49543\,
            in1 => \N__50137\,
            in2 => \N__43115\,
            in3 => \N__43067\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__46754\,
            in1 => \N__43037\,
            in2 => \_gnd_net_\,
            in3 => \N__47662\,
            lcout => \current_shift_inst.control_input_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__47661\,
            in1 => \N__46433\,
            in2 => \_gnd_net_\,
            in3 => \N__43028\,
            lcout => \current_shift_inst.control_input_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__46478\,
            in1 => \N__43016\,
            in2 => \_gnd_net_\,
            in3 => \N__47659\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__47660\,
            in1 => \_gnd_net_\,
            in2 => \N__43007\,
            in3 => \N__46448\,
            lcout => \current_shift_inst.control_input_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__50136\,
            in1 => \N__49544\,
            in2 => \N__42992\,
            in3 => \N__42947\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__42920\,
            in1 => \N__46328\,
            in2 => \_gnd_net_\,
            in3 => \N__47617\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__47618\,
            in1 => \N__46301\,
            in2 => \_gnd_net_\,
            in3 => \N__42908\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__42896\,
            in1 => \N__46271\,
            in2 => \_gnd_net_\,
            in3 => \N__47619\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__47620\,
            in1 => \N__46244\,
            in2 => \_gnd_net_\,
            in3 => \N__43187\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__43178\,
            in1 => \N__46985\,
            in2 => \_gnd_net_\,
            in3 => \N__47624\,
            lcout => \current_shift_inst.control_input_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__47623\,
            in1 => \N__43166\,
            in2 => \_gnd_net_\,
            in3 => \N__46604\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__43157\,
            in1 => \N__46184\,
            in2 => \_gnd_net_\,
            in3 => \N__47622\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__47621\,
            in1 => \N__46211\,
            in2 => \_gnd_net_\,
            in3 => \N__43148\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__47614\,
            in1 => \N__43139\,
            in2 => \_gnd_net_\,
            in3 => \N__46556\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__43127\,
            in1 => \N__46358\,
            in2 => \_gnd_net_\,
            in3 => \N__47612\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => \current_shift_inst.control_input_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43118\,
            in3 => \N__46825\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53771\,
            ce => 'H',
            sr => \N__53366\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47613\,
            lcout => \current_shift_inst.N_1619_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__47615\,
            in1 => \N__46529\,
            in2 => \_gnd_net_\,
            in3 => \N__43295\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__46502\,
            in1 => \N__47616\,
            in2 => \_gnd_net_\,
            in3 => \N__43283\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__46919\,
            in1 => \N__47665\,
            in2 => \_gnd_net_\,
            in3 => \N__43274\,
            lcout => \current_shift_inst.control_input_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__47664\,
            in1 => \N__46583\,
            in2 => \_gnd_net_\,
            in3 => \N__43262\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__47651\,
            in1 => \N__46964\,
            in2 => \_gnd_net_\,
            in3 => \N__43253\,
            lcout => \current_shift_inst.control_input_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__46661\,
            in1 => \N__43244\,
            in2 => \_gnd_net_\,
            in3 => \N__47649\,
            lcout => \current_shift_inst.control_input_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__47652\,
            in1 => \N__43235\,
            in2 => \_gnd_net_\,
            in3 => \N__46868\,
            lcout => \current_shift_inst.control_input_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__46733\,
            in1 => \N__43223\,
            in2 => \_gnd_net_\,
            in3 => \N__47648\,
            lcout => \current_shift_inst.control_input_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__47647\,
            in1 => \_gnd_net_\,
            in2 => \N__43211\,
            in3 => \N__46775\,
            lcout => \current_shift_inst.control_input_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__43199\,
            in1 => \N__46634\,
            in2 => \_gnd_net_\,
            in3 => \N__47650\,
            lcout => \current_shift_inst.control_input_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43435\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53760\,
            ce => 'H',
            sr => \N__53375\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__52236\,
            in1 => \N__47858\,
            in2 => \_gnd_net_\,
            in3 => \N__52421\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53760\,
            ce => 'H',
            sr => \N__53375\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43411\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53760\,
            ce => 'H',
            sr => \N__53375\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47698\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43381\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53749\,
            ce => 'H',
            sr => \N__53387\
        );

    \current_shift_inst.PI_CTRL.prop_term_28_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43360\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53749\,
            ce => 'H',
            sr => \N__53387\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43339\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53749\,
            ce => 'H',
            sr => \N__53387\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43309\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53749\,
            ce => 'H',
            sr => \N__53387\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__52420\,
            in1 => \N__47897\,
            in2 => \_gnd_net_\,
            in3 => \N__52238\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53749\,
            ce => 'H',
            sr => \N__53387\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43519\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53749\,
            ce => 'H',
            sr => \N__53387\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__52419\,
            in1 => \N__47918\,
            in2 => \_gnd_net_\,
            in3 => \N__52237\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53749\,
            ce => 'H',
            sr => \N__53387\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43495\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53744\,
            ce => 'H',
            sr => \N__53393\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52368\,
            in1 => \N__48047\,
            in2 => \_gnd_net_\,
            in3 => \N__52215\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53744\,
            ce => 'H',
            sr => \N__53393\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__43462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53744\,
            ce => 'H',
            sr => \N__53393\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__52371\,
            in1 => \N__52214\,
            in2 => \_gnd_net_\,
            in3 => \N__48263\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53744\,
            ce => 'H',
            sr => \N__53393\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__52211\,
            in1 => \N__52373\,
            in2 => \_gnd_net_\,
            in3 => \N__48239\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53744\,
            ce => 'H',
            sr => \N__53393\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__52369\,
            in1 => \N__52212\,
            in2 => \_gnd_net_\,
            in3 => \N__48377\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53744\,
            ce => 'H',
            sr => \N__53393\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__52210\,
            in1 => \N__52372\,
            in2 => \_gnd_net_\,
            in3 => \N__48290\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53744\,
            ce => 'H',
            sr => \N__53393\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__52370\,
            in1 => \N__52213\,
            in2 => \_gnd_net_\,
            in3 => \N__48317\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53744\,
            ce => 'H',
            sr => \N__53393\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_16_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__52204\,
            in1 => \N__52363\,
            in2 => \_gnd_net_\,
            in3 => \N__48557\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53740\,
            ce => 'H',
            sr => \N__53404\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__52206\,
            in1 => \N__52365\,
            in2 => \_gnd_net_\,
            in3 => \N__48485\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53740\,
            ce => 'H',
            sr => \N__53404\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__52362\,
            in1 => \N__52209\,
            in2 => \_gnd_net_\,
            in3 => \N__48512\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53740\,
            ce => 'H',
            sr => \N__53404\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__52207\,
            in1 => \N__52366\,
            in2 => \_gnd_net_\,
            in3 => \N__48461\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53740\,
            ce => 'H',
            sr => \N__53404\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__52361\,
            in1 => \N__52208\,
            in2 => \_gnd_net_\,
            in3 => \N__48215\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53740\,
            ce => 'H',
            sr => \N__53404\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_16_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__52205\,
            in1 => \N__52364\,
            in2 => \_gnd_net_\,
            in3 => \N__48536\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53740\,
            ce => 'H',
            sr => \N__53404\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_16_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__50950\,
            in1 => \N__51231\,
            in2 => \N__50848\,
            in3 => \N__50786\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_16_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__51230\,
            in1 => \N__50840\,
            in2 => \N__50793\,
            in3 => \N__50949\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_16_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__51140\,
            in1 => \N__51188\,
            in2 => \N__50681\,
            in3 => \N__51062\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_16_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__52187\,
            in1 => \N__52401\,
            in2 => \_gnd_net_\,
            in3 => \N__48077\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53731\,
            ce => 'H',
            sr => \N__53412\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_16_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52400\,
            in1 => \N__48104\,
            in2 => \_gnd_net_\,
            in3 => \N__52188\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53731\,
            ce => 'H',
            sr => \N__53412\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44149\,
            in2 => \N__44093\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_17_3_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__53855\,
            ce => \N__44194\,
            sr => \N__53312\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44545\,
            in2 => \N__44123\,
            in3 => \N__43658\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__53855\,
            ce => \N__44194\,
            sr => \N__53312\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44092\,
            in2 => \N__44521\,
            in3 => \N__43637\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__53855\,
            ce => \N__44194\,
            sr => \N__53312\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44546\,
            in2 => \N__44491\,
            in3 => \N__43616\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__53855\,
            ce => \N__44194\,
            sr => \N__53312\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44458\,
            in2 => \N__44522\,
            in3 => \N__43586\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__53855\,
            ce => \N__44194\,
            sr => \N__53312\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44428\,
            in2 => \N__44492\,
            in3 => \N__43559\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__53855\,
            ce => \N__44194\,
            sr => \N__53312\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44395\,
            in2 => \N__44462\,
            in3 => \N__43529\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__53855\,
            ce => \N__44194\,
            sr => \N__53312\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44362\,
            in2 => \N__44432\,
            in3 => \N__43868\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__53855\,
            ce => \N__44194\,
            sr => \N__53312\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44338\,
            in2 => \N__44402\,
            in3 => \N__43847\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_17_4_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__53854\,
            ce => \N__44195\,
            sr => \N__53313\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44314\,
            in2 => \N__44369\,
            in3 => \N__43826\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__53854\,
            ce => \N__44195\,
            sr => \N__53313\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44339\,
            in2 => \N__44776\,
            in3 => \N__43805\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__53854\,
            ce => \N__44195\,
            sr => \N__53313\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44315\,
            in2 => \N__44746\,
            in3 => \N__43784\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__53854\,
            ce => \N__44195\,
            sr => \N__53313\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44713\,
            in2 => \N__44777\,
            in3 => \N__43763\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__53854\,
            ce => \N__44195\,
            sr => \N__53313\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44686\,
            in2 => \N__44747\,
            in3 => \N__43745\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__53854\,
            ce => \N__44195\,
            sr => \N__53313\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44656\,
            in2 => \N__44717\,
            in3 => \N__43721\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__53854\,
            ce => \N__44195\,
            sr => \N__53313\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44687\,
            in2 => \N__44626\,
            in3 => \N__43697\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__53854\,
            ce => \N__44195\,
            sr => \N__53313\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44593\,
            in2 => \N__44663\,
            in3 => \N__44045\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_17_5_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__53853\,
            ce => \N__44193\,
            sr => \N__53315\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44569\,
            in2 => \N__44630\,
            in3 => \N__44024\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__53853\,
            ce => \N__44193\,
            sr => \N__53315\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44594\,
            in2 => \N__45013\,
            in3 => \N__44003\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__53853\,
            ce => \N__44193\,
            sr => \N__53315\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44570\,
            in2 => \N__44986\,
            in3 => \N__43982\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__53853\,
            ce => \N__44193\,
            sr => \N__53315\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44956\,
            in2 => \N__45014\,
            in3 => \N__43958\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__53853\,
            ce => \N__44193\,
            sr => \N__53315\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44929\,
            in2 => \N__44987\,
            in3 => \N__43937\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__53853\,
            ce => \N__44193\,
            sr => \N__53315\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44899\,
            in2 => \N__44960\,
            in3 => \N__43913\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__53853\,
            ce => \N__44193\,
            sr => \N__53315\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44866\,
            in2 => \N__44933\,
            in3 => \N__43892\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__53853\,
            ce => \N__44193\,
            sr => \N__53315\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44839\,
            in2 => \N__44906\,
            in3 => \N__44273\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_17_6_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__53850\,
            ce => \N__44182\,
            sr => \N__53316\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44818\,
            in2 => \N__44873\,
            in3 => \N__44252\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__53850\,
            ce => \N__44182\,
            sr => \N__53316\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44840\,
            in2 => \N__44798\,
            in3 => \N__44237\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__53850\,
            ce => \N__44182\,
            sr => \N__53316\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44819\,
            in2 => \N__45287\,
            in3 => \N__44219\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__53850\,
            ce => \N__44182\,
            sr => \N__53316\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44216\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53850\,
            ce => \N__44182\,
            sr => \N__53316\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45395\,
            in1 => \N__44142\,
            in2 => \_gnd_net_\,
            in3 => \N__44126\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_7_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__53846\,
            ce => \N__45268\,
            sr => \N__53317\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45390\,
            in1 => \N__44115\,
            in2 => \_gnd_net_\,
            in3 => \N__44096\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__53846\,
            ce => \N__45268\,
            sr => \N__53317\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45396\,
            in1 => \N__44082\,
            in2 => \_gnd_net_\,
            in3 => \N__44066\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__53846\,
            ce => \N__45268\,
            sr => \N__53317\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45391\,
            in1 => \N__44539\,
            in2 => \_gnd_net_\,
            in3 => \N__44525\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__53846\,
            ce => \N__45268\,
            sr => \N__53317\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45397\,
            in1 => \N__44509\,
            in2 => \_gnd_net_\,
            in3 => \N__44495\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__53846\,
            ce => \N__45268\,
            sr => \N__53317\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45392\,
            in1 => \N__44479\,
            in2 => \_gnd_net_\,
            in3 => \N__44465\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__53846\,
            ce => \N__45268\,
            sr => \N__53317\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45394\,
            in1 => \N__44451\,
            in2 => \_gnd_net_\,
            in3 => \N__44435\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__53846\,
            ce => \N__45268\,
            sr => \N__53317\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45393\,
            in1 => \N__44421\,
            in2 => \_gnd_net_\,
            in3 => \N__44405\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__53846\,
            ce => \N__45268\,
            sr => \N__53317\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45381\,
            in1 => \N__44394\,
            in2 => \_gnd_net_\,
            in3 => \N__44372\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__53841\,
            ce => \N__45251\,
            sr => \N__53318\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45407\,
            in1 => \N__44361\,
            in2 => \_gnd_net_\,
            in3 => \N__44342\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__53841\,
            ce => \N__45251\,
            sr => \N__53318\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45378\,
            in1 => \N__44332\,
            in2 => \_gnd_net_\,
            in3 => \N__44318\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__53841\,
            ce => \N__45251\,
            sr => \N__53318\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45404\,
            in1 => \N__44308\,
            in2 => \_gnd_net_\,
            in3 => \N__44294\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__53841\,
            ce => \N__45251\,
            sr => \N__53318\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45379\,
            in1 => \N__44764\,
            in2 => \_gnd_net_\,
            in3 => \N__44750\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__53841\,
            ce => \N__45251\,
            sr => \N__53318\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45405\,
            in1 => \N__44734\,
            in2 => \_gnd_net_\,
            in3 => \N__44720\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__53841\,
            ce => \N__45251\,
            sr => \N__53318\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45380\,
            in1 => \N__44706\,
            in2 => \_gnd_net_\,
            in3 => \N__44690\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__53841\,
            ce => \N__45251\,
            sr => \N__53318\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45406\,
            in1 => \N__44680\,
            in2 => \_gnd_net_\,
            in3 => \N__44666\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__53841\,
            ce => \N__45251\,
            sr => \N__53318\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45382\,
            in1 => \N__44655\,
            in2 => \_gnd_net_\,
            in3 => \N__44633\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__53834\,
            ce => \N__45269\,
            sr => \N__53320\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45386\,
            in1 => \N__44619\,
            in2 => \_gnd_net_\,
            in3 => \N__44597\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__53834\,
            ce => \N__45269\,
            sr => \N__53320\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45383\,
            in1 => \N__44587\,
            in2 => \_gnd_net_\,
            in3 => \N__44573\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__53834\,
            ce => \N__45269\,
            sr => \N__53320\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45387\,
            in1 => \N__44563\,
            in2 => \_gnd_net_\,
            in3 => \N__44549\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__53834\,
            ce => \N__45269\,
            sr => \N__53320\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45384\,
            in1 => \N__45006\,
            in2 => \_gnd_net_\,
            in3 => \N__44990\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__53834\,
            ce => \N__45269\,
            sr => \N__53320\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45388\,
            in1 => \N__44979\,
            in2 => \_gnd_net_\,
            in3 => \N__44963\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__53834\,
            ce => \N__45269\,
            sr => \N__53320\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45385\,
            in1 => \N__44955\,
            in2 => \_gnd_net_\,
            in3 => \N__44936\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__53834\,
            ce => \N__45269\,
            sr => \N__53320\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45389\,
            in1 => \N__44928\,
            in2 => \_gnd_net_\,
            in3 => \N__44909\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__53834\,
            ce => \N__45269\,
            sr => \N__53320\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45398\,
            in1 => \N__44898\,
            in2 => \_gnd_net_\,
            in3 => \N__44876\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__53829\,
            ce => \N__45267\,
            sr => \N__53322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45402\,
            in1 => \N__44865\,
            in2 => \_gnd_net_\,
            in3 => \N__44843\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__53829\,
            ce => \N__45267\,
            sr => \N__53322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45399\,
            in1 => \N__44838\,
            in2 => \_gnd_net_\,
            in3 => \N__44822\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__53829\,
            ce => \N__45267\,
            sr => \N__53322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45403\,
            in1 => \N__44817\,
            in2 => \_gnd_net_\,
            in3 => \N__44801\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__53829\,
            ce => \N__45267\,
            sr => \N__53322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45400\,
            in1 => \N__44794\,
            in2 => \_gnd_net_\,
            in3 => \N__44780\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__53829\,
            ce => \N__45267\,
            sr => \N__53322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__45283\,
            in1 => \N__45401\,
            in2 => \_gnd_net_\,
            in3 => \N__45290\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53829\,
            ce => \N__45267\,
            sr => \N__53322\
        );

    \current_shift_inst.timer_s1.counter_0_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48769\,
            in1 => \N__45216\,
            in2 => \_gnd_net_\,
            in3 => \N__45194\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__53823\,
            ce => \N__48824\,
            sr => \N__53324\
        );

    \current_shift_inst.timer_s1.counter_1_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48765\,
            in1 => \N__45180\,
            in2 => \_gnd_net_\,
            in3 => \N__45155\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__53823\,
            ce => \N__48824\,
            sr => \N__53324\
        );

    \current_shift_inst.timer_s1.counter_2_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48770\,
            in1 => \N__45145\,
            in2 => \_gnd_net_\,
            in3 => \N__45131\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__53823\,
            ce => \N__48824\,
            sr => \N__53324\
        );

    \current_shift_inst.timer_s1.counter_3_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48766\,
            in1 => \N__45121\,
            in2 => \_gnd_net_\,
            in3 => \N__45107\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__53823\,
            ce => \N__48824\,
            sr => \N__53324\
        );

    \current_shift_inst.timer_s1.counter_4_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48771\,
            in1 => \N__45091\,
            in2 => \_gnd_net_\,
            in3 => \N__45077\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__53823\,
            ce => \N__48824\,
            sr => \N__53324\
        );

    \current_shift_inst.timer_s1.counter_5_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48767\,
            in1 => \N__45061\,
            in2 => \_gnd_net_\,
            in3 => \N__45047\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__53823\,
            ce => \N__48824\,
            sr => \N__53324\
        );

    \current_shift_inst.timer_s1.counter_6_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48772\,
            in1 => \N__45033\,
            in2 => \_gnd_net_\,
            in3 => \N__45017\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__53823\,
            ce => \N__48824\,
            sr => \N__53324\
        );

    \current_shift_inst.timer_s1.counter_7_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48768\,
            in1 => \N__45637\,
            in2 => \_gnd_net_\,
            in3 => \N__45623\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__53823\,
            ce => \N__48824\,
            sr => \N__53324\
        );

    \current_shift_inst.timer_s1.counter_8_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48751\,
            in1 => \N__45615\,
            in2 => \_gnd_net_\,
            in3 => \N__45587\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__53815\,
            ce => \N__48816\,
            sr => \N__53328\
        );

    \current_shift_inst.timer_s1.counter_9_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48776\,
            in1 => \N__45570\,
            in2 => \_gnd_net_\,
            in3 => \N__45548\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__53815\,
            ce => \N__48816\,
            sr => \N__53328\
        );

    \current_shift_inst.timer_s1.counter_10_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48748\,
            in1 => \N__45534\,
            in2 => \_gnd_net_\,
            in3 => \N__45518\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__53815\,
            ce => \N__48816\,
            sr => \N__53328\
        );

    \current_shift_inst.timer_s1.counter_11_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48773\,
            in1 => \N__45508\,
            in2 => \_gnd_net_\,
            in3 => \N__45494\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__53815\,
            ce => \N__48816\,
            sr => \N__53328\
        );

    \current_shift_inst.timer_s1.counter_12_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48749\,
            in1 => \N__45484\,
            in2 => \_gnd_net_\,
            in3 => \N__45470\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__53815\,
            ce => \N__48816\,
            sr => \N__53328\
        );

    \current_shift_inst.timer_s1.counter_13_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48774\,
            in1 => \N__45454\,
            in2 => \_gnd_net_\,
            in3 => \N__45440\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__53815\,
            ce => \N__48816\,
            sr => \N__53328\
        );

    \current_shift_inst.timer_s1.counter_14_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48750\,
            in1 => \N__45424\,
            in2 => \_gnd_net_\,
            in3 => \N__45410\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__53815\,
            ce => \N__48816\,
            sr => \N__53328\
        );

    \current_shift_inst.timer_s1.counter_15_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48775\,
            in1 => \N__45904\,
            in2 => \_gnd_net_\,
            in3 => \N__45890\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__53815\,
            ce => \N__48816\,
            sr => \N__53328\
        );

    \current_shift_inst.timer_s1.counter_16_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48744\,
            in1 => \N__45882\,
            in2 => \_gnd_net_\,
            in3 => \N__45854\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__53807\,
            ce => \N__48815\,
            sr => \N__53330\
        );

    \current_shift_inst.timer_s1.counter_17_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48752\,
            in1 => \N__45843\,
            in2 => \_gnd_net_\,
            in3 => \N__45815\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__53807\,
            ce => \N__48815\,
            sr => \N__53330\
        );

    \current_shift_inst.timer_s1.counter_18_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48745\,
            in1 => \N__45801\,
            in2 => \_gnd_net_\,
            in3 => \N__45785\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__53807\,
            ce => \N__48815\,
            sr => \N__53330\
        );

    \current_shift_inst.timer_s1.counter_19_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48753\,
            in1 => \N__45775\,
            in2 => \_gnd_net_\,
            in3 => \N__45761\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__53807\,
            ce => \N__48815\,
            sr => \N__53330\
        );

    \current_shift_inst.timer_s1.counter_20_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48746\,
            in1 => \N__45747\,
            in2 => \_gnd_net_\,
            in3 => \N__45731\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__53807\,
            ce => \N__48815\,
            sr => \N__53330\
        );

    \current_shift_inst.timer_s1.counter_21_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48754\,
            in1 => \N__45715\,
            in2 => \_gnd_net_\,
            in3 => \N__45701\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__53807\,
            ce => \N__48815\,
            sr => \N__53330\
        );

    \current_shift_inst.timer_s1.counter_22_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48747\,
            in1 => \N__45687\,
            in2 => \_gnd_net_\,
            in3 => \N__45671\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__53807\,
            ce => \N__48815\,
            sr => \N__53330\
        );

    \current_shift_inst.timer_s1.counter_23_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48755\,
            in1 => \N__45661\,
            in2 => \_gnd_net_\,
            in3 => \N__45647\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__53807\,
            ce => \N__48815\,
            sr => \N__53330\
        );

    \current_shift_inst.timer_s1.counter_24_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48720\,
            in1 => \N__46158\,
            in2 => \_gnd_net_\,
            in3 => \N__46136\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__53800\,
            ce => \N__48817\,
            sr => \N__53336\
        );

    \current_shift_inst.timer_s1.counter_25_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48724\,
            in1 => \N__46125\,
            in2 => \_gnd_net_\,
            in3 => \N__46097\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__53800\,
            ce => \N__48817\,
            sr => \N__53336\
        );

    \current_shift_inst.timer_s1.counter_26_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48721\,
            in1 => \N__46087\,
            in2 => \_gnd_net_\,
            in3 => \N__46073\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__53800\,
            ce => \N__48817\,
            sr => \N__53336\
        );

    \current_shift_inst.timer_s1.counter_27_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48725\,
            in1 => \N__46063\,
            in2 => \_gnd_net_\,
            in3 => \N__46049\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__53800\,
            ce => \N__48817\,
            sr => \N__53336\
        );

    \current_shift_inst.timer_s1.counter_28_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48722\,
            in1 => \N__46036\,
            in2 => \_gnd_net_\,
            in3 => \N__46022\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__53800\,
            ce => \N__48817\,
            sr => \N__53336\
        );

    \current_shift_inst.timer_s1.counter_29_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__46009\,
            in1 => \N__48723\,
            in2 => \_gnd_net_\,
            in3 => \N__46019\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53800\,
            ce => \N__48817\,
            sr => \N__53336\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45995\,
            in2 => \N__45979\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45930\,
            in2 => \N__45959\,
            in3 => \N__46425\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46426\,
            in1 => \N__49314\,
            in2 => \N__46376\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50171\,
            in2 => \N__49499\,
            in3 => \N__46346\,
            lcout => \current_shift_inst.un38_control_input_0_s0_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49318\,
            in2 => \N__46343\,
            in3 => \N__46316\,
            lcout => \current_shift_inst.un38_control_input_0_s0_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46313\,
            in2 => \N__49500\,
            in3 => \N__46289\,
            lcout => \current_shift_inst.un38_control_input_0_s0_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49322\,
            in2 => \N__46286\,
            in3 => \N__46259\,
            lcout => \current_shift_inst.un38_control_input_0_s0_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46256\,
            in2 => \N__49501\,
            in3 => \N__46232\,
            lcout => \current_shift_inst.un38_control_input_0_s0_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49342\,
            in2 => \N__46229\,
            in3 => \N__46199\,
            lcout => \current_shift_inst.un38_control_input_0_s0_8\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46196\,
            in2 => \N__49506\,
            in3 => \N__46172\,
            lcout => \current_shift_inst.un38_control_input_0_s0_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49346\,
            in2 => \N__46619\,
            in3 => \N__46595\,
            lcout => \current_shift_inst.un38_control_input_0_s0_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46592\,
            in2 => \N__49507\,
            in3 => \N__46571\,
            lcout => \current_shift_inst.un38_control_input_0_s0_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49350\,
            in2 => \N__46568\,
            in3 => \N__46544\,
            lcout => \current_shift_inst.un38_control_input_0_s0_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46541\,
            in2 => \N__49508\,
            in3 => \N__46517\,
            lcout => \current_shift_inst.un38_control_input_0_s0_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49354\,
            in2 => \N__46514\,
            in3 => \N__46490\,
            lcout => \current_shift_inst.un38_control_input_0_s0_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46487\,
            in2 => \N__49509\,
            in3 => \N__46469\,
            lcout => \current_shift_inst.un38_control_input_0_s0_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49510\,
            in2 => \N__46466\,
            in3 => \N__46442\,
            lcout => \current_shift_inst.un38_control_input_0_s0_16\,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46439\,
            in2 => \N__49615\,
            in3 => \N__46793\,
            lcout => \current_shift_inst.un38_control_input_0_s0_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49514\,
            in2 => \N__46790\,
            in3 => \N__46763\,
            lcout => \current_shift_inst.un38_control_input_0_s0_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46760\,
            in2 => \N__49616\,
            in3 => \N__46748\,
            lcout => \current_shift_inst.un38_control_input_0_s0_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49518\,
            in2 => \N__46745\,
            in3 => \N__46718\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46715\,
            in2 => \N__49617\,
            in3 => \N__46700\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49522\,
            in2 => \N__46697\,
            in3 => \N__46676\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46673\,
            in2 => \N__49618\,
            in3 => \N__46649\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49526\,
            in2 => \N__46646\,
            in3 => \N__46622\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46997\,
            in2 => \N__49619\,
            in3 => \N__46979\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49530\,
            in2 => \N__46976\,
            in3 => \N__46952\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46949\,
            in2 => \N__49620\,
            in3 => \N__46937\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49534\,
            in2 => \N__46934\,
            in3 => \N__46910\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46907\,
            in2 => \N__49621\,
            in3 => \N__46886\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49538\,
            in2 => \N__46883\,
            in3 => \N__46859\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__46856\,
            in1 => \N__46844\,
            in2 => \N__47687\,
            in3 => \N__46835\,
            lcout => \current_shift_inst.control_input_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46832\,
            in2 => \N__46826\,
            in3 => \N__46824\,
            lcout => \current_shift_inst.control_input_1\,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47165\,
            in2 => \_gnd_net_\,
            in3 => \N__47147\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47144\,
            in2 => \_gnd_net_\,
            in3 => \N__47126\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47123\,
            in2 => \_gnd_net_\,
            in3 => \N__47105\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47102\,
            in2 => \_gnd_net_\,
            in3 => \N__47084\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47081\,
            in2 => \_gnd_net_\,
            in3 => \N__47063\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47060\,
            in2 => \_gnd_net_\,
            in3 => \N__47042\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47039\,
            in2 => \_gnd_net_\,
            in3 => \N__47021\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47018\,
            in2 => \_gnd_net_\,
            in3 => \N__47000\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47345\,
            in2 => \_gnd_net_\,
            in3 => \N__47327\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47324\,
            in2 => \_gnd_net_\,
            in3 => \N__47306\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47303\,
            in2 => \_gnd_net_\,
            in3 => \N__47285\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47282\,
            in2 => \_gnd_net_\,
            in3 => \N__47261\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47258\,
            in2 => \_gnd_net_\,
            in3 => \N__47237\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_12\,
            carryout => \current_shift_inst.control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47234\,
            in2 => \_gnd_net_\,
            in3 => \N__47213\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_13\,
            carryout => \current_shift_inst.control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47210\,
            in2 => \_gnd_net_\,
            in3 => \N__47192\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_14\,
            carryout => \current_shift_inst.control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47189\,
            in2 => \_gnd_net_\,
            in3 => \N__47168\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_21_0_\,
            carryout => \current_shift_inst.control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47519\,
            in2 => \_gnd_net_\,
            in3 => \N__47501\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_16\,
            carryout => \current_shift_inst.control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47498\,
            in2 => \_gnd_net_\,
            in3 => \N__47474\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_17\,
            carryout => \current_shift_inst.control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47471\,
            in2 => \_gnd_net_\,
            in3 => \N__47447\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_18\,
            carryout => \current_shift_inst.control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47444\,
            in2 => \_gnd_net_\,
            in3 => \N__47426\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_19\,
            carryout => \current_shift_inst.control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47423\,
            in2 => \_gnd_net_\,
            in3 => \N__47405\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_20\,
            carryout => \current_shift_inst.control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47402\,
            in2 => \_gnd_net_\,
            in3 => \N__47381\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_21\,
            carryout => \current_shift_inst.control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47378\,
            in2 => \_gnd_net_\,
            in3 => \N__47360\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_22\,
            carryout => \current_shift_inst.control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47357\,
            in2 => \_gnd_net_\,
            in3 => \N__47819\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_22_0_\,
            carryout => \current_shift_inst.control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47816\,
            in2 => \_gnd_net_\,
            in3 => \N__47798\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_24\,
            carryout => \current_shift_inst.control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47795\,
            in2 => \_gnd_net_\,
            in3 => \N__47771\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_25\,
            carryout => \current_shift_inst.control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47768\,
            in2 => \_gnd_net_\,
            in3 => \N__47750\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_26\,
            carryout => \current_shift_inst.control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47747\,
            in2 => \_gnd_net_\,
            in3 => \N__47726\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_27\,
            carryout => \current_shift_inst.control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47543\,
            in2 => \_gnd_net_\,
            in3 => \N__47711\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_28\,
            carryout => \current_shift_inst.control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__47686\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47708\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47685\,
            lcout => \current_shift_inst.control_input_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51518\,
            in2 => \N__47537\,
            in3 => \N__52223\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \bfn_17_23_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \N__53761\,
            ce => 'H',
            sr => \N__53376\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__52222\,
            in1 => \N__51555\,
            in2 => \N__47996\,
            in3 => \N__47978\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \N__53761\,
            ce => 'H',
            sr => \N__53376\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__52235\,
            in1 => \N__51618\,
            in2 => \N__47975\,
            in3 => \N__47957\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \N__53761\,
            ce => 'H',
            sr => \N__53376\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51595\,
            in2 => \N__47954\,
            in3 => \N__47936\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51771\,
            in2 => \N__47933\,
            in3 => \N__47912\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51804\,
            in2 => \N__47909\,
            in3 => \N__47891\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51315\,
            in2 => \N__47888\,
            in3 => \N__47873\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51474\,
            in2 => \N__47870\,
            in3 => \N__47852\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47849\,
            in2 => \N__51280\,
            in3 => \N__47834\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_24_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50749\,
            in2 => \N__48206\,
            in3 => \N__48176\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51378\,
            in2 => \N__48173\,
            in3 => \N__48155\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50685\,
            in2 => \N__48152\,
            in3 => \N__48122\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50629\,
            in2 => \N__48119\,
            in3 => \N__48092\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50578\,
            in2 => \N__48089\,
            in3 => \N__48065\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50522\,
            in2 => \N__48062\,
            in3 => \N__48041\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52068\,
            in2 => \N__48038\,
            in3 => \N__48020\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52462\,
            in2 => \N__48017\,
            in3 => \N__47999\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_17_25_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51436\,
            in2 => \N__48416\,
            in3 => \N__48398\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51689\,
            in2 => \N__48395\,
            in3 => \N__48371\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_17_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51748\,
            in2 => \N__48368\,
            in3 => \N__48338\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50945\,
            in2 => \N__48335\,
            in3 => \N__48311\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_17_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51656\,
            in2 => \N__48308\,
            in3 => \N__48284\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_17_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50905\,
            in2 => \N__48281\,
            in3 => \N__48257\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_17_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48254\,
            in2 => \N__50844\,
            in3 => \N__48233\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_17_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48230\,
            in2 => \N__50794\,
            in3 => \N__48209\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_17_26_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_17_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51232\,
            in2 => \N__48575\,
            in3 => \N__48551\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_17_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48548\,
            in2 => \N__51196\,
            in3 => \N__48530\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48527\,
            in2 => \N__51148\,
            in3 => \N__48506\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_17_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51096\,
            in2 => \N__48503\,
            in3 => \N__48479\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_17_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48476\,
            in2 => \N__51070\,
            in3 => \N__48455\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_er_31_LC_17_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52374\,
            in1 => \N__48452\,
            in2 => \N__48437\,
            in3 => \N__48419\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53745\,
            ce => \N__52221\,
            sr => \N__53394\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_17_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__50904\,
            in1 => \N__50526\,
            in2 => \N__51100\,
            in3 => \N__50747\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_17_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__51746\,
            in1 => \N__51660\,
            in2 => \N__51707\,
            in3 => \N__52454\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_17_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__51379\,
            in1 => \N__50571\,
            in2 => \N__52073\,
            in3 => \N__50622\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_17_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__48650\,
            in1 => \N__48644\,
            in2 => \N__48638\,
            in3 => \N__48635\,
            lcout => \current_shift_inst.PI_CTRL.N_46_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_17_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__51063\,
            in1 => \N__51141\,
            in2 => \N__50692\,
            in3 => \N__51189\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_17_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51092\,
            in2 => \_gnd_net_\,
            in3 => \N__50903\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_17_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__48629\,
            in1 => \N__50527\,
            in2 => \N__48620\,
            in3 => \N__50748\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_17_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48617\,
            in1 => \N__52388\,
            in2 => \_gnd_net_\,
            in3 => \N__52189\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53733\,
            ce => 'H',
            sr => \N__53408\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_17_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__51432\,
            in1 => \N__48884\,
            in2 => \N__52418\,
            in3 => \N__48608\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_17_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__48602\,
            in1 => \N__48593\,
            in2 => \N__48587\,
            in3 => \N__51449\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_47_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_17_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__51008\,
            in1 => \N__51401\,
            in2 => \N__48584\,
            in3 => \N__48581\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0\,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_17_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52387\,
            in2 => \N__48899\,
            in3 => \N__48896\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53733\,
            ce => 'H',
            sr => \N__53408\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_17_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__50570\,
            in1 => \N__50618\,
            in2 => \N__51377\,
            in3 => \N__52058\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_tr_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48870\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48833\,
            ce => 'H',
            sr => \N__53325\
        );

    \delay_measurement_inst.stop_timer_tr_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48871\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48833\,
            ce => 'H',
            sr => \N__53325\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__48791\,
            in1 => \N__49062\,
            in2 => \_gnd_net_\,
            in3 => \N__49031\,
            lcout => \current_shift_inst.timer_s1.N_164_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_s1_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__49084\,
            in1 => \N__49144\,
            in2 => \N__49037\,
            in3 => \N__48793\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53808\,
            ce => 'H',
            sr => \N__53331\
        );

    \current_shift_inst.timer_s1.running_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__48794\,
            in1 => \N__49032\,
            in2 => \_gnd_net_\,
            in3 => \N__49063\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53808\,
            ce => 'H',
            sr => \N__53331\
        );

    \current_shift_inst.start_timer_s1_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__49083\,
            in1 => \N__48792\,
            in2 => \_gnd_net_\,
            in3 => \N__49145\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53808\,
            ce => 'H',
            sr => \N__53331\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49061\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__50082\,
            in1 => \N__49804\,
            in2 => \N__49562\,
            in3 => \N__50164\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__50165\,
            in1 => \N__50081\,
            in2 => \N__49805\,
            in3 => \N__49459\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S1_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49143\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53793\,
            ce => 'H',
            sr => \N__53338\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49064\,
            in2 => \_gnd_net_\,
            in3 => \N__49036\,
            lcout => \current_shift_inst.timer_s1.N_163_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50185\,
            in2 => \_gnd_net_\,
            in3 => \N__51534\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53781\,
            ce => 'H',
            sr => \N__53355\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48982\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53776\,
            ce => 'H',
            sr => \N__53362\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48964\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53776\,
            ce => 'H',
            sr => \N__53362\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48940\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53776\,
            ce => 'H',
            sr => \N__53362\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48919\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53776\,
            ce => 'H',
            sr => \N__53362\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50374\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53772\,
            ce => 'H',
            sr => \N__53367\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50353\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53772\,
            ce => 'H',
            sr => \N__53367\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50329\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53772\,
            ce => 'H',
            sr => \N__53367\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50302\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53772\,
            ce => 'H',
            sr => \N__53367\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50278\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53772\,
            ce => 'H',
            sr => \N__53367\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50257\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53772\,
            ce => 'H',
            sr => \N__53367\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50233\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53772\,
            ce => 'H',
            sr => \N__53367\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50206\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53772\,
            ce => 'H',
            sr => \N__53367\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50186\,
            in2 => \N__51535\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_23_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50468\,
            in2 => \N__51562\,
            in3 => \N__50462\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__53765\,
            ce => 'H',
            sr => \N__53370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51622\,
            in2 => \N__50459\,
            in3 => \N__50450\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__53765\,
            ce => 'H',
            sr => \N__53370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50447\,
            in2 => \N__51602\,
            in3 => \N__50438\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__53765\,
            ce => 'H',
            sr => \N__53370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50435\,
            in2 => \N__51785\,
            in3 => \N__50423\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__53765\,
            ce => 'H',
            sr => \N__53370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50420\,
            in2 => \N__51818\,
            in3 => \N__50411\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__53765\,
            ce => 'H',
            sr => \N__53370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50408\,
            in2 => \N__51332\,
            in3 => \N__50399\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__53765\,
            ce => 'H',
            sr => \N__53370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50396\,
            in2 => \N__51500\,
            in3 => \N__50390\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__53765\,
            ce => 'H',
            sr => \N__53370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50387\,
            in2 => \N__51281\,
            in3 => \N__50378\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_18_24_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__53762\,
            ce => 'H',
            sr => \N__53377\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50762\,
            in2 => \N__50753\,
            in3 => \N__50720\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__53762\,
            ce => 'H',
            sr => \N__53377\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50717\,
            in2 => \N__51383\,
            in3 => \N__50708\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__53762\,
            ce => 'H',
            sr => \N__53377\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50705\,
            in2 => \N__50696\,
            in3 => \N__50648\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__53762\,
            ce => 'H',
            sr => \N__53377\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50645\,
            in2 => \N__50636\,
            in3 => \N__50594\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__53762\,
            ce => 'H',
            sr => \N__53377\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50591\,
            in2 => \N__50582\,
            in3 => \N__50549\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__53762\,
            ce => 'H',
            sr => \N__53377\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50546\,
            in2 => \N__50534\,
            in3 => \N__50501\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__53762\,
            ce => 'H',
            sr => \N__53377\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50498\,
            in2 => \N__52072\,
            in3 => \N__50489\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__53762\,
            ce => 'H',
            sr => \N__53377\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50486\,
            in2 => \N__52466\,
            in3 => \N__50471\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_18_25_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__53754\,
            ce => 'H',
            sr => \N__53383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_18_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51002\,
            in2 => \N__51443\,
            in3 => \N__50993\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__53754\,
            ce => 'H',
            sr => \N__53383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50990\,
            in2 => \N__51706\,
            in3 => \N__50978\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__53754\,
            ce => 'H',
            sr => \N__53383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_18_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50975\,
            in2 => \N__51752\,
            in3 => \N__50966\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__53754\,
            ce => 'H',
            sr => \N__53383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50963\,
            in2 => \N__50954\,
            in3 => \N__50924\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__53754\,
            ce => 'H',
            sr => \N__53383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51664\,
            in2 => \N__50921\,
            in3 => \N__50909\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__53754\,
            ce => 'H',
            sr => \N__53383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_18_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50906\,
            in2 => \N__50879\,
            in3 => \N__50864\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__53754\,
            ce => 'H',
            sr => \N__53383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_18_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50861\,
            in2 => \N__50849\,
            in3 => \N__50813\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__53754\,
            ce => 'H',
            sr => \N__53383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_18_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50810\,
            in2 => \N__50801\,
            in3 => \N__50765\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_18_26_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__53750\,
            ce => 'H',
            sr => \N__53388\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_18_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51248\,
            in2 => \N__51239\,
            in3 => \N__51212\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__53750\,
            ce => 'H',
            sr => \N__53388\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_18_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51209\,
            in2 => \N__51200\,
            in3 => \N__51167\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__53750\,
            ce => 'H',
            sr => \N__53388\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_18_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51164\,
            in2 => \N__51152\,
            in3 => \N__51119\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__53750\,
            ce => 'H',
            sr => \N__53388\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_18_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51116\,
            in2 => \N__51104\,
            in3 => \N__51074\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__53750\,
            ce => 'H',
            sr => \N__53388\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_18_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51071\,
            in2 => \N__51041\,
            in3 => \N__51026\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__53750\,
            ce => 'H',
            sr => \N__53388\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_18_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__52367\,
            in1 => \N__51023\,
            in2 => \_gnd_net_\,
            in3 => \N__51014\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53750\,
            ce => 'H',
            sr => \N__53388\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_18_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__51275\,
            in1 => \N__51814\,
            in2 => \N__51331\,
            in3 => \N__51781\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_18_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__51629\,
            in1 => \N__51496\,
            in2 => \N__51011\,
            in3 => \N__51594\,
            lcout => \current_shift_inst.PI_CTRL.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_18_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__51324\,
            in1 => \N__51813\,
            in2 => \_gnd_net_\,
            in3 => \N__51780\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_18_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__51747\,
            in1 => \N__51705\,
            in2 => \N__51668\,
            in3 => \N__52455\,
            lcout => \current_shift_inst.PI_CTRL.N_46_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_18_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010011"
        )
    port map (
            in0 => \N__51628\,
            in1 => \N__51593\,
            in2 => \N__51569\,
            in3 => \N__51539\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_18_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__51276\,
            in1 => \N__51495\,
            in2 => \N__51458\,
            in3 => \N__51455\,
            lcout => \current_shift_inst.PI_CTRL.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_18_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__52375\,
            in1 => \N__51431\,
            in2 => \_gnd_net_\,
            in3 => \N__51407\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_18_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52422\,
            in1 => \N__51395\,
            in2 => \_gnd_net_\,
            in3 => \N__52190\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53734\,
            ce => 'H',
            sr => \N__53409\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__52425\,
            in1 => \N__51341\,
            in2 => \_gnd_net_\,
            in3 => \N__52234\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53777\,
            ce => 'H',
            sr => \N__53371\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__52233\,
            in1 => \N__52426\,
            in2 => \_gnd_net_\,
            in3 => \N__51293\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53777\,
            ce => 'H',
            sr => \N__53371\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_20_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51877\,
            in2 => \_gnd_net_\,
            in3 => \N__51859\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIF9C4_12_LC_20_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52009\,
            in1 => \N__52022\,
            in2 => \N__51989\,
            in3 => \N__51974\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA4C4_10_LC_20_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__52021\,
            in1 => \N__51928\,
            in2 => \N__52010\,
            in3 => \N__51949\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPCN8_12_LC_20_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__51985\,
            in1 => \N__51973\,
            in2 => \N__51962\,
            in3 => \N__51959\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIC8E4_10_LC_20_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52622\,
            in1 => \N__51953\,
            in2 => \N__51935\,
            in3 => \N__52601\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_20_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__51907\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52648\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIT7H5_18_LC_20_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__51896\,
            in1 => \N__51842\,
            in2 => \N__51911\,
            in3 => \N__51830\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIOHB4_13_LC_20_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__51908\,
            in1 => \N__51895\,
            in2 => \N__51884\,
            in3 => \N__51863\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_20_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51841\,
            in2 => \_gnd_net_\,
            in3 => \N__51829\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7TP8_19_LC_20_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52579\,
            in1 => \N__52658\,
            in2 => \N__52652\,
            in3 => \N__52649\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_20_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52637\,
            in1 => \N__52631\,
            in2 => \N__52625\,
            in3 => \N__52484\,
            lcout => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIROF4_24_LC_20_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__52531\,
            in1 => \N__52519\,
            in2 => \N__52505\,
            in3 => \N__52621\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNITQF4_19_LC_20_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__52544\,
            in1 => \N__52600\,
            in2 => \N__52559\,
            in3 => \N__52580\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI2182_27_LC_20_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52558\,
            in2 => \_gnd_net_\,
            in3 => \N__52543\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNICPJ5_24_LC_20_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52532\,
            in1 => \N__52520\,
            in2 => \N__52508\,
            in3 => \N__52504\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_20_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52424\,
            in1 => \N__52478\,
            in2 => \_gnd_net_\,
            in3 => \N__52241\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53755\,
            ce => 'H',
            sr => \N__53395\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_21_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52427\,
            in1 => \N__52253\,
            in2 => \_gnd_net_\,
            in3 => \N__52239\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53773\,
            ce => 'H',
            sr => \N__53389\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_12_LC_22_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__52901\,
            in1 => \N__52889\,
            in2 => \N__52880\,
            in3 => \N__52865\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_23_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__54085\,
            in1 => \N__53993\,
            in2 => \N__52838\,
            in3 => \N__54259\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53835\,
            ce => 'H',
            sr => \N__53343\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__52831\,
            in1 => \N__53002\,
            in2 => \N__53056\,
            in3 => \N__52802\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => \current_shift_inst.PI_CTRL.N_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__54063\,
            in1 => \N__54165\,
            in2 => \N__52841\,
            in3 => \N__54246\,
            lcout => \current_shift_inst.PI_CTRL.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52830\,
            in2 => \_gnd_net_\,
            in3 => \N__53043\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_23_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52989\,
            in1 => \N__52699\,
            in2 => \N__52805\,
            in3 => \N__53093\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_6_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52698\,
            in2 => \_gnd_net_\,
            in3 => \N__53092\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__54091\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => pwm_duty_input_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53842\,
            ce => 'H',
            sr => \N__53347\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111010"
        )
    port map (
            in0 => \N__52703\,
            in1 => \N__53992\,
            in2 => \N__54260\,
            in3 => \N__54092\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53842\,
            ce => 'H',
            sr => \N__53347\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_24_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100100010"
        )
    port map (
            in0 => \N__54261\,
            in1 => \N__54089\,
            in2 => \N__53994\,
            in3 => \N__53091\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53836\,
            ce => 'H',
            sr => \N__53356\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_24_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__54088\,
            in1 => \N__53982\,
            in2 => \N__53057\,
            in3 => \N__54263\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53836\,
            ce => 'H',
            sr => \N__53356\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_24_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100100010"
        )
    port map (
            in0 => \N__54262\,
            in1 => \N__54090\,
            in2 => \N__53995\,
            in3 => \N__53003\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53836\,
            ce => 'H',
            sr => \N__53356\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__54116\,
            in1 => \N__53915\,
            in2 => \_gnd_net_\,
            in3 => \N__54191\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53836\,
            ce => 'H',
            sr => \N__53356\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53900\,
            in2 => \_gnd_net_\,
            in3 => \N__54177\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53836\,
            ce => 'H',
            sr => \N__53356\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_24_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010101010101"
        )
    port map (
            in0 => \N__52907\,
            in1 => \N__54167\,
            in2 => \N__53996\,
            in3 => \N__54014\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53836\,
            ce => 'H',
            sr => \N__53356\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_24_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52946\,
            in2 => \_gnd_net_\,
            in3 => \N__54178\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53836\,
            ce => 'H',
            sr => \N__53356\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_24_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__54179\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52928\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53836\,
            ce => 'H',
            sr => \N__53356\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__54166\,
            in1 => \N__54087\,
            in2 => \N__54278\,
            in3 => \N__54248\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_24_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__54274\,
            in1 => \N__54086\,
            in2 => \_gnd_net_\,
            in3 => \N__54247\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_97_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__54115\,
            in1 => \N__53911\,
            in2 => \N__54194\,
            in3 => \N__54190\,
            lcout => \current_shift_inst.PI_CTRL.N_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54164\,
            in2 => \_gnd_net_\,
            in3 => \N__54114\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_24_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__54067\,
            in1 => \N__54010\,
            in2 => \N__53999\,
            in3 => \N__53965\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53861\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53816\,
            ce => 'H',
            sr => \N__53372\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53890\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53816\,
            ce => 'H',
            sr => \N__53372\
        );
end \INTERFACE\;
