-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 12 2024 23:00:57

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    test : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    clock_output : out std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    test22 : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__51011\ : std_logic;
signal \N__51010\ : std_logic;
signal \N__51009\ : std_logic;
signal \N__51000\ : std_logic;
signal \N__50999\ : std_logic;
signal \N__50998\ : std_logic;
signal \N__50991\ : std_logic;
signal \N__50990\ : std_logic;
signal \N__50989\ : std_logic;
signal \N__50982\ : std_logic;
signal \N__50981\ : std_logic;
signal \N__50980\ : std_logic;
signal \N__50973\ : std_logic;
signal \N__50972\ : std_logic;
signal \N__50971\ : std_logic;
signal \N__50964\ : std_logic;
signal \N__50963\ : std_logic;
signal \N__50962\ : std_logic;
signal \N__50955\ : std_logic;
signal \N__50954\ : std_logic;
signal \N__50953\ : std_logic;
signal \N__50946\ : std_logic;
signal \N__50945\ : std_logic;
signal \N__50944\ : std_logic;
signal \N__50937\ : std_logic;
signal \N__50936\ : std_logic;
signal \N__50935\ : std_logic;
signal \N__50928\ : std_logic;
signal \N__50927\ : std_logic;
signal \N__50926\ : std_logic;
signal \N__50919\ : std_logic;
signal \N__50918\ : std_logic;
signal \N__50917\ : std_logic;
signal \N__50910\ : std_logic;
signal \N__50909\ : std_logic;
signal \N__50908\ : std_logic;
signal \N__50901\ : std_logic;
signal \N__50900\ : std_logic;
signal \N__50899\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50891\ : std_logic;
signal \N__50890\ : std_logic;
signal \N__50883\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50881\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50873\ : std_logic;
signal \N__50872\ : std_logic;
signal \N__50855\ : std_logic;
signal \N__50852\ : std_logic;
signal \N__50851\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50847\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50836\ : std_logic;
signal \N__50831\ : std_logic;
signal \N__50828\ : std_logic;
signal \N__50827\ : std_logic;
signal \N__50824\ : std_logic;
signal \N__50821\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50815\ : std_logic;
signal \N__50812\ : std_logic;
signal \N__50809\ : std_logic;
signal \N__50804\ : std_logic;
signal \N__50801\ : std_logic;
signal \N__50800\ : std_logic;
signal \N__50797\ : std_logic;
signal \N__50794\ : std_logic;
signal \N__50791\ : std_logic;
signal \N__50786\ : std_logic;
signal \N__50783\ : std_logic;
signal \N__50782\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50780\ : std_logic;
signal \N__50779\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50777\ : std_logic;
signal \N__50776\ : std_logic;
signal \N__50775\ : std_logic;
signal \N__50774\ : std_logic;
signal \N__50773\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50771\ : std_logic;
signal \N__50770\ : std_logic;
signal \N__50769\ : std_logic;
signal \N__50768\ : std_logic;
signal \N__50767\ : std_logic;
signal \N__50766\ : std_logic;
signal \N__50765\ : std_logic;
signal \N__50764\ : std_logic;
signal \N__50763\ : std_logic;
signal \N__50762\ : std_logic;
signal \N__50761\ : std_logic;
signal \N__50760\ : std_logic;
signal \N__50759\ : std_logic;
signal \N__50758\ : std_logic;
signal \N__50757\ : std_logic;
signal \N__50756\ : std_logic;
signal \N__50755\ : std_logic;
signal \N__50754\ : std_logic;
signal \N__50745\ : std_logic;
signal \N__50736\ : std_logic;
signal \N__50731\ : std_logic;
signal \N__50722\ : std_logic;
signal \N__50713\ : std_logic;
signal \N__50704\ : std_logic;
signal \N__50695\ : std_logic;
signal \N__50686\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50668\ : std_logic;
signal \N__50665\ : std_logic;
signal \N__50660\ : std_logic;
signal \N__50657\ : std_logic;
signal \N__50656\ : std_logic;
signal \N__50653\ : std_logic;
signal \N__50650\ : std_logic;
signal \N__50647\ : std_logic;
signal \N__50642\ : std_logic;
signal \N__50641\ : std_logic;
signal \N__50640\ : std_logic;
signal \N__50637\ : std_logic;
signal \N__50634\ : std_logic;
signal \N__50633\ : std_logic;
signal \N__50630\ : std_logic;
signal \N__50625\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50619\ : std_logic;
signal \N__50616\ : std_logic;
signal \N__50613\ : std_logic;
signal \N__50610\ : std_logic;
signal \N__50607\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50597\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50591\ : std_logic;
signal \N__50590\ : std_logic;
signal \N__50589\ : std_logic;
signal \N__50588\ : std_logic;
signal \N__50585\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50577\ : std_logic;
signal \N__50574\ : std_logic;
signal \N__50571\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50563\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50557\ : std_logic;
signal \N__50556\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50550\ : std_logic;
signal \N__50547\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50528\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50522\ : std_logic;
signal \N__50521\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50519\ : std_logic;
signal \N__50518\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50516\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50513\ : std_logic;
signal \N__50512\ : std_logic;
signal \N__50511\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50508\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50497\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50494\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50486\ : std_logic;
signal \N__50485\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50483\ : std_logic;
signal \N__50482\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50479\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50469\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50461\ : std_logic;
signal \N__50458\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50442\ : std_logic;
signal \N__50435\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50406\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50401\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50399\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50397\ : std_logic;
signal \N__50396\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50367\ : std_logic;
signal \N__50364\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50352\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50332\ : std_logic;
signal \N__50331\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50328\ : std_logic;
signal \N__50327\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50319\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50297\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50295\ : std_logic;
signal \N__50294\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50283\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50210\ : std_logic;
signal \N__50207\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50189\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50173\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50130\ : std_logic;
signal \N__50123\ : std_logic;
signal \N__50116\ : std_logic;
signal \N__50111\ : std_logic;
signal \N__50104\ : std_logic;
signal \N__50075\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50071\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50063\ : std_logic;
signal \N__50060\ : std_logic;
signal \N__50057\ : std_logic;
signal \N__50054\ : std_logic;
signal \N__50051\ : std_logic;
signal \N__50050\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50046\ : std_logic;
signal \N__50045\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50043\ : std_logic;
signal \N__50042\ : std_logic;
signal \N__50041\ : std_logic;
signal \N__50040\ : std_logic;
signal \N__50039\ : std_logic;
signal \N__50038\ : std_logic;
signal \N__50037\ : std_logic;
signal \N__50036\ : std_logic;
signal \N__50035\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50032\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50030\ : std_logic;
signal \N__50029\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50027\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50025\ : std_logic;
signal \N__50024\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50022\ : std_logic;
signal \N__50021\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50018\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50015\ : std_logic;
signal \N__50014\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50012\ : std_logic;
signal \N__50011\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50009\ : std_logic;
signal \N__50008\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50003\ : std_logic;
signal \N__50002\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49997\ : std_logic;
signal \N__49996\ : std_logic;
signal \N__49995\ : std_logic;
signal \N__49994\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49992\ : std_logic;
signal \N__49991\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49989\ : std_logic;
signal \N__49988\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49985\ : std_logic;
signal \N__49984\ : std_logic;
signal \N__49983\ : std_logic;
signal \N__49982\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49980\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49977\ : std_logic;
signal \N__49976\ : std_logic;
signal \N__49975\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49973\ : std_logic;
signal \N__49972\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49970\ : std_logic;
signal \N__49969\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49966\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49963\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49961\ : std_logic;
signal \N__49960\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49958\ : std_logic;
signal \N__49957\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49954\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49951\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49945\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49938\ : std_logic;
signal \N__49937\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49935\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49932\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49927\ : std_logic;
signal \N__49926\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49917\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49915\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49913\ : std_logic;
signal \N__49912\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49909\ : std_logic;
signal \N__49908\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49906\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49904\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49901\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49895\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49579\ : std_logic;
signal \N__49578\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49563\ : std_logic;
signal \N__49560\ : std_logic;
signal \N__49557\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49550\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49544\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49529\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49520\ : std_logic;
signal \N__49517\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49511\ : std_logic;
signal \N__49508\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49502\ : std_logic;
signal \N__49501\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49472\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49466\ : std_logic;
signal \N__49465\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49463\ : std_logic;
signal \N__49462\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49448\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49440\ : std_logic;
signal \N__49437\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49430\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49388\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49358\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49347\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49339\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49316\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49271\ : std_logic;
signal \N__49270\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49268\ : std_logic;
signal \N__49265\ : std_logic;
signal \N__49262\ : std_logic;
signal \N__49259\ : std_logic;
signal \N__49256\ : std_logic;
signal \N__49253\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49247\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49245\ : std_logic;
signal \N__49244\ : std_logic;
signal \N__49241\ : std_logic;
signal \N__49240\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49238\ : std_logic;
signal \N__49237\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49235\ : std_logic;
signal \N__49234\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49232\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49229\ : std_logic;
signal \N__49228\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49226\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49223\ : std_logic;
signal \N__49222\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49220\ : std_logic;
signal \N__49219\ : std_logic;
signal \N__49218\ : std_logic;
signal \N__49217\ : std_logic;
signal \N__49216\ : std_logic;
signal \N__49215\ : std_logic;
signal \N__49214\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49211\ : std_logic;
signal \N__49210\ : std_logic;
signal \N__49209\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49207\ : std_logic;
signal \N__49206\ : std_logic;
signal \N__49205\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49201\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49199\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49196\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49193\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49190\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49185\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49183\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49181\ : std_logic;
signal \N__49180\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49178\ : std_logic;
signal \N__49177\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49175\ : std_logic;
signal \N__49174\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49172\ : std_logic;
signal \N__49171\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49169\ : std_logic;
signal \N__49168\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49166\ : std_logic;
signal \N__49165\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49163\ : std_logic;
signal \N__49162\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49160\ : std_logic;
signal \N__49159\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49157\ : std_logic;
signal \N__49156\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49154\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49151\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49149\ : std_logic;
signal \N__49148\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49142\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49139\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49134\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49127\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49121\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49118\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49109\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49106\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49098\ : std_logic;
signal \N__49097\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49093\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49089\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48761\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48740\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48732\ : std_logic;
signal \N__48727\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48675\ : std_logic;
signal \N__48672\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48627\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48605\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48601\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48581\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48521\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48508\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48488\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48473\ : std_logic;
signal \N__48470\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48443\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48428\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48424\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48382\ : std_logic;
signal \N__48379\ : std_logic;
signal \N__48376\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48359\ : std_logic;
signal \N__48356\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48337\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48319\ : std_logic;
signal \N__48316\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48175\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48082\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48076\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48062\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48055\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47972\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47965\ : std_logic;
signal \N__47962\ : std_logic;
signal \N__47959\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47955\ : std_logic;
signal \N__47952\ : std_logic;
signal \N__47949\ : std_logic;
signal \N__47946\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47942\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47920\ : std_logic;
signal \N__47917\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47856\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47748\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47739\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47667\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47592\ : std_logic;
signal \N__47589\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47574\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47568\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47558\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47551\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47513\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47503\ : std_logic;
signal \N__47500\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47494\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47219\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47186\ : std_logic;
signal \N__47183\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47129\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47105\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47095\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47079\ : std_logic;
signal \N__47076\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47020\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46952\ : std_logic;
signal \N__46949\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46722\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46711\ : std_logic;
signal \N__46708\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46636\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46592\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46451\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46430\ : std_logic;
signal \N__46427\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46337\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46313\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46260\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46006\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45985\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45966\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45918\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45835\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45832\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45826\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45763\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45679\ : std_logic;
signal \N__45676\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45521\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45518\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45368\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45331\ : std_logic;
signal \N__45328\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45319\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45192\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45179\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45062\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44814\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44810\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44747\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44541\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44516\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44467\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44192\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44101\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44041\ : std_logic;
signal \N__44038\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44011\ : std_logic;
signal \N__44008\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43906\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43867\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43786\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43624\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43618\ : std_logic;
signal \N__43615\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43551\ : std_logic;
signal \N__43548\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43503\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43476\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43443\ : std_logic;
signal \N__43440\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43404\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43288\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43077\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43058\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42596\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42557\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42553\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42541\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42520\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42497\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42394\ : std_logic;
signal \N__42389\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42355\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42178\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42107\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42059\ : std_logic;
signal \N__42056\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41930\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41870\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41687\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41681\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41459\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41421\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41411\ : std_logic;
signal \N__41408\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41300\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41273\ : std_logic;
signal \N__41270\ : std_logic;
signal \N__41267\ : std_logic;
signal \N__41264\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40927\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40695\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40646\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40602\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40286\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39956\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39871\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39329\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39299\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39194\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38963\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38225\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_16\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_23\ : std_logic;
signal \bfn_1_20_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_1_21_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81_cascade_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_8\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_7\ : std_logic;
signal \bfn_1_22_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\ : std_logic;
signal \bfn_1_23_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\ : std_logic;
signal \bfn_1_24_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\ : std_logic;
signal \N_86_i_i\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_0\ : std_logic;
signal \bfn_2_21_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_8\ : std_logic;
signal \bfn_2_22_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_2_23_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17\ : std_logic;
signal un7_start_stop : std_logic;
signal \pwm_generator_inst.threshold_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_3_16_0_\ : std_logic;
signal \pwm_generator_inst.un14_counter_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.threshold_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.threshold_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_6\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_3_17_0_\ : std_logic;
signal \pwm_generator_inst.threshold_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96_cascade_\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \current_shift_inst.PI_CTRL.N_94\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal pwm_duty_input_7 : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \bfn_4_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_77\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal pwm_duty_input_1 : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_16\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_24\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \bfn_5_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \bfn_5_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \bfn_5_21_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \bfn_5_22_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal pwm_duty_input_8 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_158\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\ : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_160\ : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt18\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNIDC91B_0_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt30\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal s3_phy_c : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt18\ : std_logic;
signal \bfn_10_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_start_g\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.test_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_inst2.N_58\ : std_logic;
signal \phase_controller_inst2.N_51_0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal s4_phy_c : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \elapsed_time_ns_1_RNIED91B_0_2\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.N_49_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal start_stop_c : std_logic;
signal il_max_comp2_c : std_logic;
signal \phase_controller_inst1_N_54_cascade_\ : std_logic;
signal \phase_controller_inst2.N_54\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_166_i\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \current_shift_inst.control_input_axb_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_16\ : std_logic;
signal \bfn_11_21_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_24\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_31\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal test22_c : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14\ : std_logic;
signal \phase_controller_inst1.N_52\ : std_logic;
signal \phase_controller_inst1_N_54\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.N_1271_i\ : std_logic;
signal \current_shift_inst.control_input_1\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\ : std_logic;
signal \current_shift_inst.control_input_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\ : std_logic;
signal \current_shift_inst.control_input_cry_14\ : std_logic;
signal \current_shift_inst.control_input_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\ : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\ : std_logic;
signal \current_shift_inst.control_input_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\ : std_logic;
signal \current_shift_inst.control_input_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\ : std_logic;
signal \current_shift_inst.control_input_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\ : std_logic;
signal \current_shift_inst.control_input_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\ : std_logic;
signal \current_shift_inst.control_input_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\ : std_logic;
signal \current_shift_inst.control_input_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\ : std_logic;
signal \current_shift_inst.control_input_cry_22\ : std_logic;
signal \current_shift_inst.control_input_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\ : std_logic;
signal \current_shift_inst.control_input_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\ : std_logic;
signal \current_shift_inst.control_input_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\ : std_logic;
signal \current_shift_inst.control_input_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\ : std_logic;
signal \current_shift_inst.control_input_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\ : std_logic;
signal \current_shift_inst.control_input_cry_28\ : std_logic;
signal \current_shift_inst.control_input_cry_29\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\ : std_logic;
signal \pll_inst.red_c_i\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \phase_controller_inst1.N_56\ : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\ : std_logic;
signal \phase_controller_inst1.test_0_sqmuxa\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_165_i\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal il_max_comp1_c : std_logic;
signal test_c : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \current_shift_inst.control_input_axb_16\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \current_shift_inst.control_input_axb_18\ : std_logic;
signal \current_shift_inst.control_input_axb_17\ : std_logic;
signal \current_shift_inst.control_input_axb_20\ : std_logic;
signal \current_shift_inst.control_input_axb_21\ : std_logic;
signal \current_shift_inst.control_input_axb_22\ : std_logic;
signal \current_shift_inst.control_input_axb_27\ : std_logic;
signal \current_shift_inst.control_input_axb_26\ : std_logic;
signal \current_shift_inst.control_input_axb_25\ : std_logic;
signal \current_shift_inst.control_input_axb_29\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal s1_phy_c : std_logic;
signal state_3 : std_logic;
signal \current_shift_inst.timer_s1.N_161_i\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_14_4_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_16\ : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt18\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_8\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_axb_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.control_input_axb_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_15_5_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_15_6_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt18\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_8\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_15\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_14\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.control_input_axb_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_16\ : std_logic;
signal \current_shift_inst.control_input_axb_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_17\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_17\ : std_logic;
signal \current_shift_inst.control_input_axb_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_18\ : std_logic;
signal \current_shift_inst.control_input_axb_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.control_input_axb_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30\ : std_logic;
signal \elapsed_time_ns_1_RNIE03T9_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt28\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \bfn_16_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \bfn_16_20_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_164_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \bfn_18_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \bfn_18_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \bfn_18_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \bfn_18_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_163_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \elapsed_time_ns_1_RNIDV2T9_0_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_start_g\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \bfn_18_21_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \bfn_18_22_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.N_161_i_g\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_18_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_18_24_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_18_25_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_18_26_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_162_i\ : std_logic;
signal \GB_BUFFER_clock_output_0_THRU_CO\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clock_output_0 : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal clock_output_wire : std_logic;
signal test_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal test22_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    clock_output <= clock_output_wire;
    test <= test_wire;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    test22 <= test22_wire;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ <= \N__30764\&\N__30791\&\N__30821\&\N__30848\&\N__30881\&\N__30911\&\N__30941\&\N__30971\&\N__30512\&\N__30542\&\N__30569\&\N__30599\&\N__30632\&\N__30662\&\N__30698\&\N__30728\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__44834\&'0'&\N__44833\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__20333\&\N__20326\&\N__20331\&\N__20325\&\N__20332\&\N__20324\&\N__20334\&\N__20321\&\N__20327\&\N__20320\&\N__20328\&\N__20322\&\N__20329\&\N__20323\&\N__20330\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__44964\&\N__44894\&'0'&'0'&'0'&\N__44892\&\N__44963\&\N__44893\&\N__44962\;
    \pwm_generator_inst.un2_threshold_2_1_16\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_2_1_15\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_2_14\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_2_13\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ <= '0'&\N__20343\&\N__20362\&\N__20344\&\N__20363\&\N__20345\&\N__25107\&\N__25319\&\N__22061\&\N__21845\&\N__21718\&\N__21792\&\N__21746\&\N__26026\&\N__22559\&\N__22589\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__44714\&\N__44711\&'0'&'0'&'0'&\N__44709\&\N__44713\&\N__44710\&\N__44712\;
    \pwm_generator_inst.un2_threshold_1_25\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_1_24\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_1_23\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_1_22\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_1_21\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_1_20\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(0);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ <= '0'&\N__30242\&\N__30275\&\N__30299\&\N__30329\&\N__30359\&\N__30389\&\N__30422\&\N__30448\&\N__30488\&\N__30071\&\N__30107\&\N__30137\&\N__30170\&\N__30206\&\N__29636\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__44815\&'0'&\N__44814\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(19);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(18);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(17);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(16);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.un1_integrator\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__27917\,
            RESETB => \N__33224\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clock_output_0
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__44835\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__44832\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__44965\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__44891\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__44715\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__44708\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__44816\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__44813\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__51009\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51011\,
            DIN => \N__51010\,
            DOUT => \N__51009\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__51011\,
            PADOUT => \N__51010\,
            PADIN => \N__51009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clock_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51000\,
            DIN => \N__50999\,
            DOUT => \N__50998\,
            PACKAGEPIN => clock_output_wire
        );

    \clock_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51000\,
            PADOUT => \N__50999\,
            PADIN => \N__50998\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__50597\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \test_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50991\,
            DIN => \N__50990\,
            DOUT => \N__50989\,
            PACKAGEPIN => test_wire
        );

    \test_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50991\,
            PADOUT => \N__50990\,
            PADIN => \N__50989\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35621\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50982\,
            DIN => \N__50981\,
            DOUT => \N__50980\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50982\,
            PADOUT => \N__50981\,
            PADIN => \N__50980\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50973\,
            DIN => \N__50972\,
            DOUT => \N__50971\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50973\,
            PADOUT => \N__50972\,
            PADIN => \N__50971\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50964\,
            DIN => \N__50963\,
            DOUT => \N__50962\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50964\,
            PADOUT => \N__50963\,
            PADIN => \N__50962\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21620\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50955\,
            DIN => \N__50954\,
            DOUT => \N__50953\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50955\,
            PADOUT => \N__50954\,
            PADIN => \N__50953\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50946\,
            DIN => \N__50945\,
            DOUT => \N__50944\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50946\,
            PADOUT => \N__50945\,
            PADIN => \N__50944\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35774\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \test22_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50937\,
            DIN => \N__50936\,
            DOUT => \N__50935\,
            PACKAGEPIN => test22_wire
        );

    \test22_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50937\,
            PADOUT => \N__50936\,
            PADIN => \N__50935\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31007\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50928\,
            DIN => \N__50927\,
            DOUT => \N__50926\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50928\,
            PADOUT => \N__50927\,
            PADIN => \N__50926\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50919\,
            DIN => \N__50918\,
            DOUT => \N__50917\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50919\,
            PADOUT => \N__50918\,
            PADIN => \N__50917\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35924\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50910\,
            DIN => \N__50909\,
            DOUT => \N__50908\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50910\,
            PADOUT => \N__50909\,
            PADIN => \N__50908\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28994\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50901\,
            DIN => \N__50900\,
            DOUT => \N__50899\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50901\,
            PADOUT => \N__50900\,
            PADIN => \N__50899\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50892\,
            DIN => \N__50891\,
            DOUT => \N__50890\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50892\,
            PADOUT => \N__50891\,
            PADIN => \N__50890\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27938\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50883\,
            DIN => \N__50882\,
            DOUT => \N__50881\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50883\,
            PADOUT => \N__50882\,
            PADIN => \N__50881\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50874\,
            DIN => \N__50873\,
            DOUT => \N__50872\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50874\,
            PADOUT => \N__50873\,
            PADIN => \N__50872\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__12164\ : CascadeMux
    port map (
            O => \N__50855\,
            I => \N__50852\
        );

    \I__12163\ : InMux
    port map (
            O => \N__50852\,
            I => \N__50847\
        );

    \I__12162\ : InMux
    port map (
            O => \N__50851\,
            I => \N__50844\
        );

    \I__12161\ : InMux
    port map (
            O => \N__50850\,
            I => \N__50841\
        );

    \I__12160\ : LocalMux
    port map (
            O => \N__50847\,
            I => \N__50836\
        );

    \I__12159\ : LocalMux
    port map (
            O => \N__50844\,
            I => \N__50836\
        );

    \I__12158\ : LocalMux
    port map (
            O => \N__50841\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__12157\ : Odrv12
    port map (
            O => \N__50836\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__12156\ : InMux
    port map (
            O => \N__50831\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__12155\ : CascadeMux
    port map (
            O => \N__50828\,
            I => \N__50824\
        );

    \I__12154\ : CascadeMux
    port map (
            O => \N__50827\,
            I => \N__50821\
        );

    \I__12153\ : InMux
    port map (
            O => \N__50824\,
            I => \N__50815\
        );

    \I__12152\ : InMux
    port map (
            O => \N__50821\,
            I => \N__50815\
        );

    \I__12151\ : InMux
    port map (
            O => \N__50820\,
            I => \N__50812\
        );

    \I__12150\ : LocalMux
    port map (
            O => \N__50815\,
            I => \N__50809\
        );

    \I__12149\ : LocalMux
    port map (
            O => \N__50812\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__12148\ : Odrv12
    port map (
            O => \N__50809\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__12147\ : InMux
    port map (
            O => \N__50804\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__12146\ : InMux
    port map (
            O => \N__50801\,
            I => \N__50797\
        );

    \I__12145\ : InMux
    port map (
            O => \N__50800\,
            I => \N__50794\
        );

    \I__12144\ : LocalMux
    port map (
            O => \N__50797\,
            I => \N__50791\
        );

    \I__12143\ : LocalMux
    port map (
            O => \N__50794\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__12142\ : Odrv12
    port map (
            O => \N__50791\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__12141\ : InMux
    port map (
            O => \N__50786\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__12140\ : InMux
    port map (
            O => \N__50783\,
            I => \N__50745\
        );

    \I__12139\ : InMux
    port map (
            O => \N__50782\,
            I => \N__50745\
        );

    \I__12138\ : InMux
    port map (
            O => \N__50781\,
            I => \N__50745\
        );

    \I__12137\ : InMux
    port map (
            O => \N__50780\,
            I => \N__50745\
        );

    \I__12136\ : InMux
    port map (
            O => \N__50779\,
            I => \N__50736\
        );

    \I__12135\ : InMux
    port map (
            O => \N__50778\,
            I => \N__50736\
        );

    \I__12134\ : InMux
    port map (
            O => \N__50777\,
            I => \N__50736\
        );

    \I__12133\ : InMux
    port map (
            O => \N__50776\,
            I => \N__50736\
        );

    \I__12132\ : InMux
    port map (
            O => \N__50775\,
            I => \N__50731\
        );

    \I__12131\ : InMux
    port map (
            O => \N__50774\,
            I => \N__50731\
        );

    \I__12130\ : InMux
    port map (
            O => \N__50773\,
            I => \N__50722\
        );

    \I__12129\ : InMux
    port map (
            O => \N__50772\,
            I => \N__50722\
        );

    \I__12128\ : InMux
    port map (
            O => \N__50771\,
            I => \N__50722\
        );

    \I__12127\ : InMux
    port map (
            O => \N__50770\,
            I => \N__50722\
        );

    \I__12126\ : InMux
    port map (
            O => \N__50769\,
            I => \N__50713\
        );

    \I__12125\ : InMux
    port map (
            O => \N__50768\,
            I => \N__50713\
        );

    \I__12124\ : InMux
    port map (
            O => \N__50767\,
            I => \N__50713\
        );

    \I__12123\ : InMux
    port map (
            O => \N__50766\,
            I => \N__50713\
        );

    \I__12122\ : InMux
    port map (
            O => \N__50765\,
            I => \N__50704\
        );

    \I__12121\ : InMux
    port map (
            O => \N__50764\,
            I => \N__50704\
        );

    \I__12120\ : InMux
    port map (
            O => \N__50763\,
            I => \N__50704\
        );

    \I__12119\ : InMux
    port map (
            O => \N__50762\,
            I => \N__50704\
        );

    \I__12118\ : InMux
    port map (
            O => \N__50761\,
            I => \N__50695\
        );

    \I__12117\ : InMux
    port map (
            O => \N__50760\,
            I => \N__50695\
        );

    \I__12116\ : InMux
    port map (
            O => \N__50759\,
            I => \N__50695\
        );

    \I__12115\ : InMux
    port map (
            O => \N__50758\,
            I => \N__50695\
        );

    \I__12114\ : InMux
    port map (
            O => \N__50757\,
            I => \N__50686\
        );

    \I__12113\ : InMux
    port map (
            O => \N__50756\,
            I => \N__50686\
        );

    \I__12112\ : InMux
    port map (
            O => \N__50755\,
            I => \N__50686\
        );

    \I__12111\ : InMux
    port map (
            O => \N__50754\,
            I => \N__50686\
        );

    \I__12110\ : LocalMux
    port map (
            O => \N__50745\,
            I => \N__50673\
        );

    \I__12109\ : LocalMux
    port map (
            O => \N__50736\,
            I => \N__50673\
        );

    \I__12108\ : LocalMux
    port map (
            O => \N__50731\,
            I => \N__50673\
        );

    \I__12107\ : LocalMux
    port map (
            O => \N__50722\,
            I => \N__50673\
        );

    \I__12106\ : LocalMux
    port map (
            O => \N__50713\,
            I => \N__50673\
        );

    \I__12105\ : LocalMux
    port map (
            O => \N__50704\,
            I => \N__50673\
        );

    \I__12104\ : LocalMux
    port map (
            O => \N__50695\,
            I => \N__50668\
        );

    \I__12103\ : LocalMux
    port map (
            O => \N__50686\,
            I => \N__50668\
        );

    \I__12102\ : Span4Mux_v
    port map (
            O => \N__50673\,
            I => \N__50665\
        );

    \I__12101\ : Odrv12
    port map (
            O => \N__50668\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__12100\ : Odrv4
    port map (
            O => \N__50665\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__12099\ : InMux
    port map (
            O => \N__50660\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__12098\ : InMux
    port map (
            O => \N__50657\,
            I => \N__50653\
        );

    \I__12097\ : InMux
    port map (
            O => \N__50656\,
            I => \N__50650\
        );

    \I__12096\ : LocalMux
    port map (
            O => \N__50653\,
            I => \N__50647\
        );

    \I__12095\ : LocalMux
    port map (
            O => \N__50650\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__12094\ : Odrv12
    port map (
            O => \N__50647\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__12093\ : CEMux
    port map (
            O => \N__50642\,
            I => \N__50637\
        );

    \I__12092\ : CEMux
    port map (
            O => \N__50641\,
            I => \N__50634\
        );

    \I__12091\ : CEMux
    port map (
            O => \N__50640\,
            I => \N__50630\
        );

    \I__12090\ : LocalMux
    port map (
            O => \N__50637\,
            I => \N__50625\
        );

    \I__12089\ : LocalMux
    port map (
            O => \N__50634\,
            I => \N__50625\
        );

    \I__12088\ : CEMux
    port map (
            O => \N__50633\,
            I => \N__50622\
        );

    \I__12087\ : LocalMux
    port map (
            O => \N__50630\,
            I => \N__50619\
        );

    \I__12086\ : Span4Mux_v
    port map (
            O => \N__50625\,
            I => \N__50616\
        );

    \I__12085\ : LocalMux
    port map (
            O => \N__50622\,
            I => \N__50613\
        );

    \I__12084\ : Span4Mux_h
    port map (
            O => \N__50619\,
            I => \N__50610\
        );

    \I__12083\ : Span4Mux_h
    port map (
            O => \N__50616\,
            I => \N__50607\
        );

    \I__12082\ : Span4Mux_h
    port map (
            O => \N__50613\,
            I => \N__50604\
        );

    \I__12081\ : Odrv4
    port map (
            O => \N__50610\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__12080\ : Odrv4
    port map (
            O => \N__50607\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__12079\ : Odrv4
    port map (
            O => \N__50604\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__12078\ : IoInMux
    port map (
            O => \N__50597\,
            I => \N__50594\
        );

    \I__12077\ : LocalMux
    port map (
            O => \N__50594\,
            I => \GB_BUFFER_clock_output_0_THRU_CO\
        );

    \I__12076\ : InMux
    port map (
            O => \N__50591\,
            I => \N__50585\
        );

    \I__12075\ : InMux
    port map (
            O => \N__50590\,
            I => \N__50580\
        );

    \I__12074\ : InMux
    port map (
            O => \N__50589\,
            I => \N__50580\
        );

    \I__12073\ : InMux
    port map (
            O => \N__50588\,
            I => \N__50577\
        );

    \I__12072\ : LocalMux
    port map (
            O => \N__50585\,
            I => \N__50574\
        );

    \I__12071\ : LocalMux
    port map (
            O => \N__50580\,
            I => \N__50571\
        );

    \I__12070\ : LocalMux
    port map (
            O => \N__50577\,
            I => \N__50568\
        );

    \I__12069\ : Span4Mux_v
    port map (
            O => \N__50574\,
            I => \N__50563\
        );

    \I__12068\ : Span4Mux_v
    port map (
            O => \N__50571\,
            I => \N__50563\
        );

    \I__12067\ : Odrv4
    port map (
            O => \N__50568\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__12066\ : Odrv4
    port map (
            O => \N__50563\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__12065\ : InMux
    port map (
            O => \N__50558\,
            I => \N__50553\
        );

    \I__12064\ : InMux
    port map (
            O => \N__50557\,
            I => \N__50550\
        );

    \I__12063\ : InMux
    port map (
            O => \N__50556\,
            I => \N__50547\
        );

    \I__12062\ : LocalMux
    port map (
            O => \N__50553\,
            I => \N__50544\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__50550\,
            I => \N__50541\
        );

    \I__12060\ : LocalMux
    port map (
            O => \N__50547\,
            I => \N__50536\
        );

    \I__12059\ : Span4Mux_v
    port map (
            O => \N__50544\,
            I => \N__50536\
        );

    \I__12058\ : Span12Mux_s9_h
    port map (
            O => \N__50541\,
            I => \N__50533\
        );

    \I__12057\ : Odrv4
    port map (
            O => \N__50536\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__12056\ : Odrv12
    port map (
            O => \N__50533\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__12055\ : InMux
    port map (
            O => \N__50528\,
            I => \N__50502\
        );

    \I__12054\ : InMux
    port map (
            O => \N__50527\,
            I => \N__50490\
        );

    \I__12053\ : InMux
    port map (
            O => \N__50526\,
            I => \N__50487\
        );

    \I__12052\ : CascadeMux
    port map (
            O => \N__50525\,
            I => \N__50474\
        );

    \I__12051\ : InMux
    port map (
            O => \N__50524\,
            I => \N__50470\
        );

    \I__12050\ : InMux
    port map (
            O => \N__50523\,
            I => \N__50464\
        );

    \I__12049\ : InMux
    port map (
            O => \N__50522\,
            I => \N__50464\
        );

    \I__12048\ : InMux
    port map (
            O => \N__50521\,
            I => \N__50461\
        );

    \I__12047\ : InMux
    port map (
            O => \N__50520\,
            I => \N__50458\
        );

    \I__12046\ : InMux
    port map (
            O => \N__50519\,
            I => \N__50449\
        );

    \I__12045\ : InMux
    port map (
            O => \N__50518\,
            I => \N__50449\
        );

    \I__12044\ : InMux
    port map (
            O => \N__50517\,
            I => \N__50449\
        );

    \I__12043\ : InMux
    port map (
            O => \N__50516\,
            I => \N__50449\
        );

    \I__12042\ : InMux
    port map (
            O => \N__50515\,
            I => \N__50442\
        );

    \I__12041\ : InMux
    port map (
            O => \N__50514\,
            I => \N__50442\
        );

    \I__12040\ : InMux
    port map (
            O => \N__50513\,
            I => \N__50442\
        );

    \I__12039\ : InMux
    port map (
            O => \N__50512\,
            I => \N__50435\
        );

    \I__12038\ : InMux
    port map (
            O => \N__50511\,
            I => \N__50435\
        );

    \I__12037\ : InMux
    port map (
            O => \N__50510\,
            I => \N__50435\
        );

    \I__12036\ : InMux
    port map (
            O => \N__50509\,
            I => \N__50424\
        );

    \I__12035\ : InMux
    port map (
            O => \N__50508\,
            I => \N__50424\
        );

    \I__12034\ : InMux
    port map (
            O => \N__50507\,
            I => \N__50424\
        );

    \I__12033\ : InMux
    port map (
            O => \N__50506\,
            I => \N__50424\
        );

    \I__12032\ : InMux
    port map (
            O => \N__50505\,
            I => \N__50424\
        );

    \I__12031\ : LocalMux
    port map (
            O => \N__50502\,
            I => \N__50421\
        );

    \I__12030\ : InMux
    port map (
            O => \N__50501\,
            I => \N__50417\
        );

    \I__12029\ : InMux
    port map (
            O => \N__50500\,
            I => \N__50412\
        );

    \I__12028\ : InMux
    port map (
            O => \N__50499\,
            I => \N__50412\
        );

    \I__12027\ : CascadeMux
    port map (
            O => \N__50498\,
            I => \N__50391\
        );

    \I__12026\ : InMux
    port map (
            O => \N__50497\,
            I => \N__50381\
        );

    \I__12025\ : InMux
    port map (
            O => \N__50496\,
            I => \N__50381\
        );

    \I__12024\ : InMux
    port map (
            O => \N__50495\,
            I => \N__50381\
        );

    \I__12023\ : InMux
    port map (
            O => \N__50494\,
            I => \N__50381\
        );

    \I__12022\ : InMux
    port map (
            O => \N__50493\,
            I => \N__50378\
        );

    \I__12021\ : LocalMux
    port map (
            O => \N__50490\,
            I => \N__50375\
        );

    \I__12020\ : LocalMux
    port map (
            O => \N__50487\,
            I => \N__50372\
        );

    \I__12019\ : InMux
    port map (
            O => \N__50486\,
            I => \N__50367\
        );

    \I__12018\ : InMux
    port map (
            O => \N__50485\,
            I => \N__50367\
        );

    \I__12017\ : InMux
    port map (
            O => \N__50484\,
            I => \N__50364\
        );

    \I__12016\ : InMux
    port map (
            O => \N__50483\,
            I => \N__50355\
        );

    \I__12015\ : InMux
    port map (
            O => \N__50482\,
            I => \N__50355\
        );

    \I__12014\ : InMux
    port map (
            O => \N__50481\,
            I => \N__50355\
        );

    \I__12013\ : InMux
    port map (
            O => \N__50480\,
            I => \N__50355\
        );

    \I__12012\ : InMux
    port map (
            O => \N__50479\,
            I => \N__50340\
        );

    \I__12011\ : InMux
    port map (
            O => \N__50478\,
            I => \N__50340\
        );

    \I__12010\ : InMux
    port map (
            O => \N__50477\,
            I => \N__50340\
        );

    \I__12009\ : InMux
    port map (
            O => \N__50474\,
            I => \N__50340\
        );

    \I__12008\ : InMux
    port map (
            O => \N__50473\,
            I => \N__50340\
        );

    \I__12007\ : LocalMux
    port map (
            O => \N__50470\,
            I => \N__50337\
        );

    \I__12006\ : InMux
    port map (
            O => \N__50469\,
            I => \N__50334\
        );

    \I__12005\ : LocalMux
    port map (
            O => \N__50464\,
            I => \N__50322\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__50461\,
            I => \N__50319\
        );

    \I__12003\ : LocalMux
    port map (
            O => \N__50458\,
            I => \N__50314\
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__50449\,
            I => \N__50314\
        );

    \I__12001\ : LocalMux
    port map (
            O => \N__50442\,
            I => \N__50311\
        );

    \I__12000\ : LocalMux
    port map (
            O => \N__50435\,
            I => \N__50304\
        );

    \I__11999\ : LocalMux
    port map (
            O => \N__50424\,
            I => \N__50304\
        );

    \I__11998\ : Span4Mux_h
    port map (
            O => \N__50421\,
            I => \N__50304\
        );

    \I__11997\ : CascadeMux
    port map (
            O => \N__50420\,
            I => \N__50299\
        );

    \I__11996\ : LocalMux
    port map (
            O => \N__50417\,
            I => \N__50287\
        );

    \I__11995\ : LocalMux
    port map (
            O => \N__50412\,
            I => \N__50284\
        );

    \I__11994\ : InMux
    port map (
            O => \N__50411\,
            I => \N__50276\
        );

    \I__11993\ : InMux
    port map (
            O => \N__50410\,
            I => \N__50276\
        );

    \I__11992\ : InMux
    port map (
            O => \N__50409\,
            I => \N__50265\
        );

    \I__11991\ : InMux
    port map (
            O => \N__50408\,
            I => \N__50265\
        );

    \I__11990\ : InMux
    port map (
            O => \N__50407\,
            I => \N__50265\
        );

    \I__11989\ : InMux
    port map (
            O => \N__50406\,
            I => \N__50265\
        );

    \I__11988\ : InMux
    port map (
            O => \N__50405\,
            I => \N__50265\
        );

    \I__11987\ : InMux
    port map (
            O => \N__50404\,
            I => \N__50256\
        );

    \I__11986\ : InMux
    port map (
            O => \N__50403\,
            I => \N__50256\
        );

    \I__11985\ : InMux
    port map (
            O => \N__50402\,
            I => \N__50256\
        );

    \I__11984\ : InMux
    port map (
            O => \N__50401\,
            I => \N__50256\
        );

    \I__11983\ : InMux
    port map (
            O => \N__50400\,
            I => \N__50251\
        );

    \I__11982\ : InMux
    port map (
            O => \N__50399\,
            I => \N__50251\
        );

    \I__11981\ : InMux
    port map (
            O => \N__50398\,
            I => \N__50248\
        );

    \I__11980\ : InMux
    port map (
            O => \N__50397\,
            I => \N__50245\
        );

    \I__11979\ : InMux
    port map (
            O => \N__50396\,
            I => \N__50234\
        );

    \I__11978\ : InMux
    port map (
            O => \N__50395\,
            I => \N__50234\
        );

    \I__11977\ : InMux
    port map (
            O => \N__50394\,
            I => \N__50234\
        );

    \I__11976\ : InMux
    port map (
            O => \N__50391\,
            I => \N__50234\
        );

    \I__11975\ : InMux
    port map (
            O => \N__50390\,
            I => \N__50234\
        );

    \I__11974\ : LocalMux
    port map (
            O => \N__50381\,
            I => \N__50219\
        );

    \I__11973\ : LocalMux
    port map (
            O => \N__50378\,
            I => \N__50219\
        );

    \I__11972\ : Span4Mux_s3_v
    port map (
            O => \N__50375\,
            I => \N__50219\
        );

    \I__11971\ : Span4Mux_v
    port map (
            O => \N__50372\,
            I => \N__50219\
        );

    \I__11970\ : LocalMux
    port map (
            O => \N__50367\,
            I => \N__50219\
        );

    \I__11969\ : LocalMux
    port map (
            O => \N__50364\,
            I => \N__50219\
        );

    \I__11968\ : LocalMux
    port map (
            O => \N__50355\,
            I => \N__50219\
        );

    \I__11967\ : InMux
    port map (
            O => \N__50354\,
            I => \N__50210\
        );

    \I__11966\ : InMux
    port map (
            O => \N__50353\,
            I => \N__50210\
        );

    \I__11965\ : InMux
    port map (
            O => \N__50352\,
            I => \N__50210\
        );

    \I__11964\ : InMux
    port map (
            O => \N__50351\,
            I => \N__50210\
        );

    \I__11963\ : LocalMux
    port map (
            O => \N__50340\,
            I => \N__50207\
        );

    \I__11962\ : Span4Mux_v
    port map (
            O => \N__50337\,
            I => \N__50202\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__50334\,
            I => \N__50202\
        );

    \I__11960\ : InMux
    port map (
            O => \N__50333\,
            I => \N__50189\
        );

    \I__11959\ : InMux
    port map (
            O => \N__50332\,
            I => \N__50189\
        );

    \I__11958\ : InMux
    port map (
            O => \N__50331\,
            I => \N__50189\
        );

    \I__11957\ : InMux
    port map (
            O => \N__50330\,
            I => \N__50189\
        );

    \I__11956\ : InMux
    port map (
            O => \N__50329\,
            I => \N__50189\
        );

    \I__11955\ : InMux
    port map (
            O => \N__50328\,
            I => \N__50189\
        );

    \I__11954\ : InMux
    port map (
            O => \N__50327\,
            I => \N__50182\
        );

    \I__11953\ : InMux
    port map (
            O => \N__50326\,
            I => \N__50182\
        );

    \I__11952\ : InMux
    port map (
            O => \N__50325\,
            I => \N__50182\
        );

    \I__11951\ : Span4Mux_h
    port map (
            O => \N__50322\,
            I => \N__50173\
        );

    \I__11950\ : Span4Mux_v
    port map (
            O => \N__50319\,
            I => \N__50173\
        );

    \I__11949\ : Span4Mux_v
    port map (
            O => \N__50314\,
            I => \N__50173\
        );

    \I__11948\ : Span4Mux_v
    port map (
            O => \N__50311\,
            I => \N__50173\
        );

    \I__11947\ : Span4Mux_v
    port map (
            O => \N__50304\,
            I => \N__50170\
        );

    \I__11946\ : InMux
    port map (
            O => \N__50303\,
            I => \N__50165\
        );

    \I__11945\ : InMux
    port map (
            O => \N__50302\,
            I => \N__50165\
        );

    \I__11944\ : InMux
    port map (
            O => \N__50299\,
            I => \N__50160\
        );

    \I__11943\ : InMux
    port map (
            O => \N__50298\,
            I => \N__50160\
        );

    \I__11942\ : InMux
    port map (
            O => \N__50297\,
            I => \N__50151\
        );

    \I__11941\ : InMux
    port map (
            O => \N__50296\,
            I => \N__50151\
        );

    \I__11940\ : InMux
    port map (
            O => \N__50295\,
            I => \N__50151\
        );

    \I__11939\ : InMux
    port map (
            O => \N__50294\,
            I => \N__50151\
        );

    \I__11938\ : InMux
    port map (
            O => \N__50293\,
            I => \N__50142\
        );

    \I__11937\ : InMux
    port map (
            O => \N__50292\,
            I => \N__50142\
        );

    \I__11936\ : InMux
    port map (
            O => \N__50291\,
            I => \N__50142\
        );

    \I__11935\ : InMux
    port map (
            O => \N__50290\,
            I => \N__50142\
        );

    \I__11934\ : Span4Mux_v
    port map (
            O => \N__50287\,
            I => \N__50137\
        );

    \I__11933\ : Span4Mux_h
    port map (
            O => \N__50284\,
            I => \N__50137\
        );

    \I__11932\ : InMux
    port map (
            O => \N__50283\,
            I => \N__50130\
        );

    \I__11931\ : InMux
    port map (
            O => \N__50282\,
            I => \N__50130\
        );

    \I__11930\ : InMux
    port map (
            O => \N__50281\,
            I => \N__50130\
        );

    \I__11929\ : LocalMux
    port map (
            O => \N__50276\,
            I => \N__50123\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__50265\,
            I => \N__50123\
        );

    \I__11927\ : LocalMux
    port map (
            O => \N__50256\,
            I => \N__50123\
        );

    \I__11926\ : LocalMux
    port map (
            O => \N__50251\,
            I => \N__50116\
        );

    \I__11925\ : LocalMux
    port map (
            O => \N__50248\,
            I => \N__50116\
        );

    \I__11924\ : LocalMux
    port map (
            O => \N__50245\,
            I => \N__50116\
        );

    \I__11923\ : LocalMux
    port map (
            O => \N__50234\,
            I => \N__50111\
        );

    \I__11922\ : Span4Mux_v
    port map (
            O => \N__50219\,
            I => \N__50111\
        );

    \I__11921\ : LocalMux
    port map (
            O => \N__50210\,
            I => \N__50104\
        );

    \I__11920\ : Span4Mux_v
    port map (
            O => \N__50207\,
            I => \N__50104\
        );

    \I__11919\ : Span4Mux_h
    port map (
            O => \N__50202\,
            I => \N__50104\
        );

    \I__11918\ : LocalMux
    port map (
            O => \N__50189\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11917\ : LocalMux
    port map (
            O => \N__50182\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11916\ : Odrv4
    port map (
            O => \N__50173\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11915\ : Odrv4
    port map (
            O => \N__50170\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11914\ : LocalMux
    port map (
            O => \N__50165\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11913\ : LocalMux
    port map (
            O => \N__50160\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11912\ : LocalMux
    port map (
            O => \N__50151\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11911\ : LocalMux
    port map (
            O => \N__50142\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11910\ : Odrv4
    port map (
            O => \N__50137\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11909\ : LocalMux
    port map (
            O => \N__50130\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11908\ : Odrv4
    port map (
            O => \N__50123\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11907\ : Odrv12
    port map (
            O => \N__50116\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11906\ : Odrv4
    port map (
            O => \N__50111\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11905\ : Odrv4
    port map (
            O => \N__50104\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11904\ : CascadeMux
    port map (
            O => \N__50075\,
            I => \N__50071\
        );

    \I__11903\ : CascadeMux
    port map (
            O => \N__50074\,
            I => \N__50068\
        );

    \I__11902\ : InMux
    port map (
            O => \N__50071\,
            I => \N__50063\
        );

    \I__11901\ : InMux
    port map (
            O => \N__50068\,
            I => \N__50063\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__50063\,
            I => \N__50060\
        );

    \I__11899\ : Span4Mux_h
    port map (
            O => \N__50060\,
            I => \N__50057\
        );

    \I__11898\ : Odrv4
    port map (
            O => \N__50057\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\
        );

    \I__11897\ : InMux
    port map (
            O => \N__50054\,
            I => \N__50051\
        );

    \I__11896\ : LocalMux
    port map (
            O => \N__50051\,
            I => \N__49896\
        );

    \I__11895\ : ClkMux
    port map (
            O => \N__50050\,
            I => \N__49583\
        );

    \I__11894\ : ClkMux
    port map (
            O => \N__50049\,
            I => \N__49583\
        );

    \I__11893\ : ClkMux
    port map (
            O => \N__50048\,
            I => \N__49583\
        );

    \I__11892\ : ClkMux
    port map (
            O => \N__50047\,
            I => \N__49583\
        );

    \I__11891\ : ClkMux
    port map (
            O => \N__50046\,
            I => \N__49583\
        );

    \I__11890\ : ClkMux
    port map (
            O => \N__50045\,
            I => \N__49583\
        );

    \I__11889\ : ClkMux
    port map (
            O => \N__50044\,
            I => \N__49583\
        );

    \I__11888\ : ClkMux
    port map (
            O => \N__50043\,
            I => \N__49583\
        );

    \I__11887\ : ClkMux
    port map (
            O => \N__50042\,
            I => \N__49583\
        );

    \I__11886\ : ClkMux
    port map (
            O => \N__50041\,
            I => \N__49583\
        );

    \I__11885\ : ClkMux
    port map (
            O => \N__50040\,
            I => \N__49583\
        );

    \I__11884\ : ClkMux
    port map (
            O => \N__50039\,
            I => \N__49583\
        );

    \I__11883\ : ClkMux
    port map (
            O => \N__50038\,
            I => \N__49583\
        );

    \I__11882\ : ClkMux
    port map (
            O => \N__50037\,
            I => \N__49583\
        );

    \I__11881\ : ClkMux
    port map (
            O => \N__50036\,
            I => \N__49583\
        );

    \I__11880\ : ClkMux
    port map (
            O => \N__50035\,
            I => \N__49583\
        );

    \I__11879\ : ClkMux
    port map (
            O => \N__50034\,
            I => \N__49583\
        );

    \I__11878\ : ClkMux
    port map (
            O => \N__50033\,
            I => \N__49583\
        );

    \I__11877\ : ClkMux
    port map (
            O => \N__50032\,
            I => \N__49583\
        );

    \I__11876\ : ClkMux
    port map (
            O => \N__50031\,
            I => \N__49583\
        );

    \I__11875\ : ClkMux
    port map (
            O => \N__50030\,
            I => \N__49583\
        );

    \I__11874\ : ClkMux
    port map (
            O => \N__50029\,
            I => \N__49583\
        );

    \I__11873\ : ClkMux
    port map (
            O => \N__50028\,
            I => \N__49583\
        );

    \I__11872\ : ClkMux
    port map (
            O => \N__50027\,
            I => \N__49583\
        );

    \I__11871\ : ClkMux
    port map (
            O => \N__50026\,
            I => \N__49583\
        );

    \I__11870\ : ClkMux
    port map (
            O => \N__50025\,
            I => \N__49583\
        );

    \I__11869\ : ClkMux
    port map (
            O => \N__50024\,
            I => \N__49583\
        );

    \I__11868\ : ClkMux
    port map (
            O => \N__50023\,
            I => \N__49583\
        );

    \I__11867\ : ClkMux
    port map (
            O => \N__50022\,
            I => \N__49583\
        );

    \I__11866\ : ClkMux
    port map (
            O => \N__50021\,
            I => \N__49583\
        );

    \I__11865\ : ClkMux
    port map (
            O => \N__50020\,
            I => \N__49583\
        );

    \I__11864\ : ClkMux
    port map (
            O => \N__50019\,
            I => \N__49583\
        );

    \I__11863\ : ClkMux
    port map (
            O => \N__50018\,
            I => \N__49583\
        );

    \I__11862\ : ClkMux
    port map (
            O => \N__50017\,
            I => \N__49583\
        );

    \I__11861\ : ClkMux
    port map (
            O => \N__50016\,
            I => \N__49583\
        );

    \I__11860\ : ClkMux
    port map (
            O => \N__50015\,
            I => \N__49583\
        );

    \I__11859\ : ClkMux
    port map (
            O => \N__50014\,
            I => \N__49583\
        );

    \I__11858\ : ClkMux
    port map (
            O => \N__50013\,
            I => \N__49583\
        );

    \I__11857\ : ClkMux
    port map (
            O => \N__50012\,
            I => \N__49583\
        );

    \I__11856\ : ClkMux
    port map (
            O => \N__50011\,
            I => \N__49583\
        );

    \I__11855\ : ClkMux
    port map (
            O => \N__50010\,
            I => \N__49583\
        );

    \I__11854\ : ClkMux
    port map (
            O => \N__50009\,
            I => \N__49583\
        );

    \I__11853\ : ClkMux
    port map (
            O => \N__50008\,
            I => \N__49583\
        );

    \I__11852\ : ClkMux
    port map (
            O => \N__50007\,
            I => \N__49583\
        );

    \I__11851\ : ClkMux
    port map (
            O => \N__50006\,
            I => \N__49583\
        );

    \I__11850\ : ClkMux
    port map (
            O => \N__50005\,
            I => \N__49583\
        );

    \I__11849\ : ClkMux
    port map (
            O => \N__50004\,
            I => \N__49583\
        );

    \I__11848\ : ClkMux
    port map (
            O => \N__50003\,
            I => \N__49583\
        );

    \I__11847\ : ClkMux
    port map (
            O => \N__50002\,
            I => \N__49583\
        );

    \I__11846\ : ClkMux
    port map (
            O => \N__50001\,
            I => \N__49583\
        );

    \I__11845\ : ClkMux
    port map (
            O => \N__50000\,
            I => \N__49583\
        );

    \I__11844\ : ClkMux
    port map (
            O => \N__49999\,
            I => \N__49583\
        );

    \I__11843\ : ClkMux
    port map (
            O => \N__49998\,
            I => \N__49583\
        );

    \I__11842\ : ClkMux
    port map (
            O => \N__49997\,
            I => \N__49583\
        );

    \I__11841\ : ClkMux
    port map (
            O => \N__49996\,
            I => \N__49583\
        );

    \I__11840\ : ClkMux
    port map (
            O => \N__49995\,
            I => \N__49583\
        );

    \I__11839\ : ClkMux
    port map (
            O => \N__49994\,
            I => \N__49583\
        );

    \I__11838\ : ClkMux
    port map (
            O => \N__49993\,
            I => \N__49583\
        );

    \I__11837\ : ClkMux
    port map (
            O => \N__49992\,
            I => \N__49583\
        );

    \I__11836\ : ClkMux
    port map (
            O => \N__49991\,
            I => \N__49583\
        );

    \I__11835\ : ClkMux
    port map (
            O => \N__49990\,
            I => \N__49583\
        );

    \I__11834\ : ClkMux
    port map (
            O => \N__49989\,
            I => \N__49583\
        );

    \I__11833\ : ClkMux
    port map (
            O => \N__49988\,
            I => \N__49583\
        );

    \I__11832\ : ClkMux
    port map (
            O => \N__49987\,
            I => \N__49583\
        );

    \I__11831\ : ClkMux
    port map (
            O => \N__49986\,
            I => \N__49583\
        );

    \I__11830\ : ClkMux
    port map (
            O => \N__49985\,
            I => \N__49583\
        );

    \I__11829\ : ClkMux
    port map (
            O => \N__49984\,
            I => \N__49583\
        );

    \I__11828\ : ClkMux
    port map (
            O => \N__49983\,
            I => \N__49583\
        );

    \I__11827\ : ClkMux
    port map (
            O => \N__49982\,
            I => \N__49583\
        );

    \I__11826\ : ClkMux
    port map (
            O => \N__49981\,
            I => \N__49583\
        );

    \I__11825\ : ClkMux
    port map (
            O => \N__49980\,
            I => \N__49583\
        );

    \I__11824\ : ClkMux
    port map (
            O => \N__49979\,
            I => \N__49583\
        );

    \I__11823\ : ClkMux
    port map (
            O => \N__49978\,
            I => \N__49583\
        );

    \I__11822\ : ClkMux
    port map (
            O => \N__49977\,
            I => \N__49583\
        );

    \I__11821\ : ClkMux
    port map (
            O => \N__49976\,
            I => \N__49583\
        );

    \I__11820\ : ClkMux
    port map (
            O => \N__49975\,
            I => \N__49583\
        );

    \I__11819\ : ClkMux
    port map (
            O => \N__49974\,
            I => \N__49583\
        );

    \I__11818\ : ClkMux
    port map (
            O => \N__49973\,
            I => \N__49583\
        );

    \I__11817\ : ClkMux
    port map (
            O => \N__49972\,
            I => \N__49583\
        );

    \I__11816\ : ClkMux
    port map (
            O => \N__49971\,
            I => \N__49583\
        );

    \I__11815\ : ClkMux
    port map (
            O => \N__49970\,
            I => \N__49583\
        );

    \I__11814\ : ClkMux
    port map (
            O => \N__49969\,
            I => \N__49583\
        );

    \I__11813\ : ClkMux
    port map (
            O => \N__49968\,
            I => \N__49583\
        );

    \I__11812\ : ClkMux
    port map (
            O => \N__49967\,
            I => \N__49583\
        );

    \I__11811\ : ClkMux
    port map (
            O => \N__49966\,
            I => \N__49583\
        );

    \I__11810\ : ClkMux
    port map (
            O => \N__49965\,
            I => \N__49583\
        );

    \I__11809\ : ClkMux
    port map (
            O => \N__49964\,
            I => \N__49583\
        );

    \I__11808\ : ClkMux
    port map (
            O => \N__49963\,
            I => \N__49583\
        );

    \I__11807\ : ClkMux
    port map (
            O => \N__49962\,
            I => \N__49583\
        );

    \I__11806\ : ClkMux
    port map (
            O => \N__49961\,
            I => \N__49583\
        );

    \I__11805\ : ClkMux
    port map (
            O => \N__49960\,
            I => \N__49583\
        );

    \I__11804\ : ClkMux
    port map (
            O => \N__49959\,
            I => \N__49583\
        );

    \I__11803\ : ClkMux
    port map (
            O => \N__49958\,
            I => \N__49583\
        );

    \I__11802\ : ClkMux
    port map (
            O => \N__49957\,
            I => \N__49583\
        );

    \I__11801\ : ClkMux
    port map (
            O => \N__49956\,
            I => \N__49583\
        );

    \I__11800\ : ClkMux
    port map (
            O => \N__49955\,
            I => \N__49583\
        );

    \I__11799\ : ClkMux
    port map (
            O => \N__49954\,
            I => \N__49583\
        );

    \I__11798\ : ClkMux
    port map (
            O => \N__49953\,
            I => \N__49583\
        );

    \I__11797\ : ClkMux
    port map (
            O => \N__49952\,
            I => \N__49583\
        );

    \I__11796\ : ClkMux
    port map (
            O => \N__49951\,
            I => \N__49583\
        );

    \I__11795\ : ClkMux
    port map (
            O => \N__49950\,
            I => \N__49583\
        );

    \I__11794\ : ClkMux
    port map (
            O => \N__49949\,
            I => \N__49583\
        );

    \I__11793\ : ClkMux
    port map (
            O => \N__49948\,
            I => \N__49583\
        );

    \I__11792\ : ClkMux
    port map (
            O => \N__49947\,
            I => \N__49583\
        );

    \I__11791\ : ClkMux
    port map (
            O => \N__49946\,
            I => \N__49583\
        );

    \I__11790\ : ClkMux
    port map (
            O => \N__49945\,
            I => \N__49583\
        );

    \I__11789\ : ClkMux
    port map (
            O => \N__49944\,
            I => \N__49583\
        );

    \I__11788\ : ClkMux
    port map (
            O => \N__49943\,
            I => \N__49583\
        );

    \I__11787\ : ClkMux
    port map (
            O => \N__49942\,
            I => \N__49583\
        );

    \I__11786\ : ClkMux
    port map (
            O => \N__49941\,
            I => \N__49583\
        );

    \I__11785\ : ClkMux
    port map (
            O => \N__49940\,
            I => \N__49583\
        );

    \I__11784\ : ClkMux
    port map (
            O => \N__49939\,
            I => \N__49583\
        );

    \I__11783\ : ClkMux
    port map (
            O => \N__49938\,
            I => \N__49583\
        );

    \I__11782\ : ClkMux
    port map (
            O => \N__49937\,
            I => \N__49583\
        );

    \I__11781\ : ClkMux
    port map (
            O => \N__49936\,
            I => \N__49583\
        );

    \I__11780\ : ClkMux
    port map (
            O => \N__49935\,
            I => \N__49583\
        );

    \I__11779\ : ClkMux
    port map (
            O => \N__49934\,
            I => \N__49583\
        );

    \I__11778\ : ClkMux
    port map (
            O => \N__49933\,
            I => \N__49583\
        );

    \I__11777\ : ClkMux
    port map (
            O => \N__49932\,
            I => \N__49583\
        );

    \I__11776\ : ClkMux
    port map (
            O => \N__49931\,
            I => \N__49583\
        );

    \I__11775\ : ClkMux
    port map (
            O => \N__49930\,
            I => \N__49583\
        );

    \I__11774\ : ClkMux
    port map (
            O => \N__49929\,
            I => \N__49583\
        );

    \I__11773\ : ClkMux
    port map (
            O => \N__49928\,
            I => \N__49583\
        );

    \I__11772\ : ClkMux
    port map (
            O => \N__49927\,
            I => \N__49583\
        );

    \I__11771\ : ClkMux
    port map (
            O => \N__49926\,
            I => \N__49583\
        );

    \I__11770\ : ClkMux
    port map (
            O => \N__49925\,
            I => \N__49583\
        );

    \I__11769\ : ClkMux
    port map (
            O => \N__49924\,
            I => \N__49583\
        );

    \I__11768\ : ClkMux
    port map (
            O => \N__49923\,
            I => \N__49583\
        );

    \I__11767\ : ClkMux
    port map (
            O => \N__49922\,
            I => \N__49583\
        );

    \I__11766\ : ClkMux
    port map (
            O => \N__49921\,
            I => \N__49583\
        );

    \I__11765\ : ClkMux
    port map (
            O => \N__49920\,
            I => \N__49583\
        );

    \I__11764\ : ClkMux
    port map (
            O => \N__49919\,
            I => \N__49583\
        );

    \I__11763\ : ClkMux
    port map (
            O => \N__49918\,
            I => \N__49583\
        );

    \I__11762\ : ClkMux
    port map (
            O => \N__49917\,
            I => \N__49583\
        );

    \I__11761\ : ClkMux
    port map (
            O => \N__49916\,
            I => \N__49583\
        );

    \I__11760\ : ClkMux
    port map (
            O => \N__49915\,
            I => \N__49583\
        );

    \I__11759\ : ClkMux
    port map (
            O => \N__49914\,
            I => \N__49583\
        );

    \I__11758\ : ClkMux
    port map (
            O => \N__49913\,
            I => \N__49583\
        );

    \I__11757\ : ClkMux
    port map (
            O => \N__49912\,
            I => \N__49583\
        );

    \I__11756\ : ClkMux
    port map (
            O => \N__49911\,
            I => \N__49583\
        );

    \I__11755\ : ClkMux
    port map (
            O => \N__49910\,
            I => \N__49583\
        );

    \I__11754\ : ClkMux
    port map (
            O => \N__49909\,
            I => \N__49583\
        );

    \I__11753\ : ClkMux
    port map (
            O => \N__49908\,
            I => \N__49583\
        );

    \I__11752\ : ClkMux
    port map (
            O => \N__49907\,
            I => \N__49583\
        );

    \I__11751\ : ClkMux
    port map (
            O => \N__49906\,
            I => \N__49583\
        );

    \I__11750\ : ClkMux
    port map (
            O => \N__49905\,
            I => \N__49583\
        );

    \I__11749\ : ClkMux
    port map (
            O => \N__49904\,
            I => \N__49583\
        );

    \I__11748\ : ClkMux
    port map (
            O => \N__49903\,
            I => \N__49583\
        );

    \I__11747\ : ClkMux
    port map (
            O => \N__49902\,
            I => \N__49583\
        );

    \I__11746\ : ClkMux
    port map (
            O => \N__49901\,
            I => \N__49583\
        );

    \I__11745\ : ClkMux
    port map (
            O => \N__49900\,
            I => \N__49583\
        );

    \I__11744\ : ClkMux
    port map (
            O => \N__49899\,
            I => \N__49583\
        );

    \I__11743\ : Glb2LocalMux
    port map (
            O => \N__49896\,
            I => \N__49583\
        );

    \I__11742\ : ClkMux
    port map (
            O => \N__49895\,
            I => \N__49583\
        );

    \I__11741\ : ClkMux
    port map (
            O => \N__49894\,
            I => \N__49583\
        );

    \I__11740\ : GlobalMux
    port map (
            O => \N__49583\,
            I => clock_output_0
        );

    \I__11739\ : InMux
    port map (
            O => \N__49580\,
            I => \N__49570\
        );

    \I__11738\ : InMux
    port map (
            O => \N__49579\,
            I => \N__49570\
        );

    \I__11737\ : InMux
    port map (
            O => \N__49578\,
            I => \N__49570\
        );

    \I__11736\ : CEMux
    port map (
            O => \N__49577\,
            I => \N__49567\
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__49570\,
            I => \N__49560\
        );

    \I__11734\ : LocalMux
    port map (
            O => \N__49567\,
            I => \N__49557\
        );

    \I__11733\ : CEMux
    port map (
            O => \N__49566\,
            I => \N__49554\
        );

    \I__11732\ : CEMux
    port map (
            O => \N__49565\,
            I => \N__49551\
        );

    \I__11731\ : CEMux
    port map (
            O => \N__49564\,
            I => \N__49545\
        );

    \I__11730\ : CEMux
    port map (
            O => \N__49563\,
            I => \N__49539\
        );

    \I__11729\ : Span4Mux_v
    port map (
            O => \N__49560\,
            I => \N__49530\
        );

    \I__11728\ : Span4Mux_h
    port map (
            O => \N__49557\,
            I => \N__49530\
        );

    \I__11727\ : LocalMux
    port map (
            O => \N__49554\,
            I => \N__49530\
        );

    \I__11726\ : LocalMux
    port map (
            O => \N__49551\,
            I => \N__49530\
        );

    \I__11725\ : CEMux
    port map (
            O => \N__49550\,
            I => \N__49517\
        );

    \I__11724\ : CEMux
    port map (
            O => \N__49549\,
            I => \N__49514\
        );

    \I__11723\ : CEMux
    port map (
            O => \N__49548\,
            I => \N__49511\
        );

    \I__11722\ : LocalMux
    port map (
            O => \N__49545\,
            I => \N__49508\
        );

    \I__11721\ : CEMux
    port map (
            O => \N__49544\,
            I => \N__49505\
        );

    \I__11720\ : CEMux
    port map (
            O => \N__49543\,
            I => \N__49502\
        );

    \I__11719\ : CEMux
    port map (
            O => \N__49542\,
            I => \N__49497\
        );

    \I__11718\ : LocalMux
    port map (
            O => \N__49539\,
            I => \N__49494\
        );

    \I__11717\ : Span4Mux_v
    port map (
            O => \N__49530\,
            I => \N__49491\
        );

    \I__11716\ : InMux
    port map (
            O => \N__49529\,
            I => \N__49482\
        );

    \I__11715\ : InMux
    port map (
            O => \N__49528\,
            I => \N__49482\
        );

    \I__11714\ : InMux
    port map (
            O => \N__49527\,
            I => \N__49482\
        );

    \I__11713\ : InMux
    port map (
            O => \N__49526\,
            I => \N__49482\
        );

    \I__11712\ : InMux
    port map (
            O => \N__49525\,
            I => \N__49473\
        );

    \I__11711\ : InMux
    port map (
            O => \N__49524\,
            I => \N__49473\
        );

    \I__11710\ : InMux
    port map (
            O => \N__49523\,
            I => \N__49473\
        );

    \I__11709\ : InMux
    port map (
            O => \N__49522\,
            I => \N__49473\
        );

    \I__11708\ : CEMux
    port map (
            O => \N__49521\,
            I => \N__49466\
        );

    \I__11707\ : CEMux
    port map (
            O => \N__49520\,
            I => \N__49457\
        );

    \I__11706\ : LocalMux
    port map (
            O => \N__49517\,
            I => \N__49454\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__49514\,
            I => \N__49451\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__49511\,
            I => \N__49448\
        );

    \I__11703\ : Span4Mux_h
    port map (
            O => \N__49508\,
            I => \N__49443\
        );

    \I__11702\ : LocalMux
    port map (
            O => \N__49505\,
            I => \N__49443\
        );

    \I__11701\ : LocalMux
    port map (
            O => \N__49502\,
            I => \N__49440\
        );

    \I__11700\ : CEMux
    port map (
            O => \N__49501\,
            I => \N__49437\
        );

    \I__11699\ : CEMux
    port map (
            O => \N__49500\,
            I => \N__49430\
        );

    \I__11698\ : LocalMux
    port map (
            O => \N__49497\,
            I => \N__49426\
        );

    \I__11697\ : Span4Mux_h
    port map (
            O => \N__49494\,
            I => \N__49417\
        );

    \I__11696\ : Span4Mux_h
    port map (
            O => \N__49491\,
            I => \N__49417\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__49482\,
            I => \N__49417\
        );

    \I__11694\ : LocalMux
    port map (
            O => \N__49473\,
            I => \N__49417\
        );

    \I__11693\ : InMux
    port map (
            O => \N__49472\,
            I => \N__49408\
        );

    \I__11692\ : InMux
    port map (
            O => \N__49471\,
            I => \N__49408\
        );

    \I__11691\ : InMux
    port map (
            O => \N__49470\,
            I => \N__49408\
        );

    \I__11690\ : InMux
    port map (
            O => \N__49469\,
            I => \N__49408\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__49466\,
            I => \N__49405\
        );

    \I__11688\ : CEMux
    port map (
            O => \N__49465\,
            I => \N__49402\
        );

    \I__11687\ : InMux
    port map (
            O => \N__49464\,
            I => \N__49393\
        );

    \I__11686\ : InMux
    port map (
            O => \N__49463\,
            I => \N__49393\
        );

    \I__11685\ : InMux
    port map (
            O => \N__49462\,
            I => \N__49393\
        );

    \I__11684\ : InMux
    port map (
            O => \N__49461\,
            I => \N__49393\
        );

    \I__11683\ : CEMux
    port map (
            O => \N__49460\,
            I => \N__49390\
        );

    \I__11682\ : LocalMux
    port map (
            O => \N__49457\,
            I => \N__49378\
        );

    \I__11681\ : Span4Mux_h
    port map (
            O => \N__49454\,
            I => \N__49378\
        );

    \I__11680\ : Span4Mux_h
    port map (
            O => \N__49451\,
            I => \N__49378\
        );

    \I__11679\ : Span4Mux_h
    port map (
            O => \N__49448\,
            I => \N__49378\
        );

    \I__11678\ : Span4Mux_v
    port map (
            O => \N__49443\,
            I => \N__49375\
        );

    \I__11677\ : Span4Mux_v
    port map (
            O => \N__49440\,
            I => \N__49372\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__49437\,
            I => \N__49369\
        );

    \I__11675\ : InMux
    port map (
            O => \N__49436\,
            I => \N__49360\
        );

    \I__11674\ : InMux
    port map (
            O => \N__49435\,
            I => \N__49360\
        );

    \I__11673\ : InMux
    port map (
            O => \N__49434\,
            I => \N__49360\
        );

    \I__11672\ : InMux
    port map (
            O => \N__49433\,
            I => \N__49360\
        );

    \I__11671\ : LocalMux
    port map (
            O => \N__49430\,
            I => \N__49353\
        );

    \I__11670\ : InMux
    port map (
            O => \N__49429\,
            I => \N__49350\
        );

    \I__11669\ : Span4Mux_v
    port map (
            O => \N__49426\,
            I => \N__49347\
        );

    \I__11668\ : Span4Mux_v
    port map (
            O => \N__49417\,
            I => \N__49342\
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__49408\,
            I => \N__49342\
        );

    \I__11666\ : Span4Mux_s2_v
    port map (
            O => \N__49405\,
            I => \N__49339\
        );

    \I__11665\ : LocalMux
    port map (
            O => \N__49402\,
            I => \N__49334\
        );

    \I__11664\ : LocalMux
    port map (
            O => \N__49393\,
            I => \N__49334\
        );

    \I__11663\ : LocalMux
    port map (
            O => \N__49390\,
            I => \N__49331\
        );

    \I__11662\ : InMux
    port map (
            O => \N__49389\,
            I => \N__49324\
        );

    \I__11661\ : InMux
    port map (
            O => \N__49388\,
            I => \N__49324\
        );

    \I__11660\ : InMux
    port map (
            O => \N__49387\,
            I => \N__49324\
        );

    \I__11659\ : Span4Mux_v
    port map (
            O => \N__49378\,
            I => \N__49321\
        );

    \I__11658\ : Span4Mux_s1_v
    port map (
            O => \N__49375\,
            I => \N__49316\
        );

    \I__11657\ : Span4Mux_h
    port map (
            O => \N__49372\,
            I => \N__49316\
        );

    \I__11656\ : Span4Mux_h
    port map (
            O => \N__49369\,
            I => \N__49311\
        );

    \I__11655\ : LocalMux
    port map (
            O => \N__49360\,
            I => \N__49311\
        );

    \I__11654\ : InMux
    port map (
            O => \N__49359\,
            I => \N__49302\
        );

    \I__11653\ : InMux
    port map (
            O => \N__49358\,
            I => \N__49302\
        );

    \I__11652\ : InMux
    port map (
            O => \N__49357\,
            I => \N__49302\
        );

    \I__11651\ : InMux
    port map (
            O => \N__49356\,
            I => \N__49302\
        );

    \I__11650\ : Span4Mux_v
    port map (
            O => \N__49353\,
            I => \N__49297\
        );

    \I__11649\ : LocalMux
    port map (
            O => \N__49350\,
            I => \N__49297\
        );

    \I__11648\ : Span4Mux_h
    port map (
            O => \N__49347\,
            I => \N__49288\
        );

    \I__11647\ : Span4Mux_v
    port map (
            O => \N__49342\,
            I => \N__49288\
        );

    \I__11646\ : Span4Mux_h
    port map (
            O => \N__49339\,
            I => \N__49288\
        );

    \I__11645\ : Span4Mux_h
    port map (
            O => \N__49334\,
            I => \N__49288\
        );

    \I__11644\ : Odrv12
    port map (
            O => \N__49331\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11643\ : LocalMux
    port map (
            O => \N__49324\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11642\ : Odrv4
    port map (
            O => \N__49321\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11641\ : Odrv4
    port map (
            O => \N__49316\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11640\ : Odrv4
    port map (
            O => \N__49311\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__49302\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11638\ : Odrv4
    port map (
            O => \N__49297\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11637\ : Odrv4
    port map (
            O => \N__49288\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11636\ : InMux
    port map (
            O => \N__49271\,
            I => \N__49265\
        );

    \I__11635\ : InMux
    port map (
            O => \N__49270\,
            I => \N__49262\
        );

    \I__11634\ : InMux
    port map (
            O => \N__49269\,
            I => \N__49259\
        );

    \I__11633\ : InMux
    port map (
            O => \N__49268\,
            I => \N__49256\
        );

    \I__11632\ : LocalMux
    port map (
            O => \N__49265\,
            I => \N__49253\
        );

    \I__11631\ : LocalMux
    port map (
            O => \N__49262\,
            I => \N__49250\
        );

    \I__11630\ : LocalMux
    port map (
            O => \N__49259\,
            I => \N__49247\
        );

    \I__11629\ : LocalMux
    port map (
            O => \N__49256\,
            I => \N__49241\
        );

    \I__11628\ : Glb2LocalMux
    port map (
            O => \N__49253\,
            I => \N__48767\
        );

    \I__11627\ : Glb2LocalMux
    port map (
            O => \N__49250\,
            I => \N__48767\
        );

    \I__11626\ : Glb2LocalMux
    port map (
            O => \N__49247\,
            I => \N__48767\
        );

    \I__11625\ : SRMux
    port map (
            O => \N__49246\,
            I => \N__48767\
        );

    \I__11624\ : SRMux
    port map (
            O => \N__49245\,
            I => \N__48767\
        );

    \I__11623\ : SRMux
    port map (
            O => \N__49244\,
            I => \N__48767\
        );

    \I__11622\ : Glb2LocalMux
    port map (
            O => \N__49241\,
            I => \N__48767\
        );

    \I__11621\ : SRMux
    port map (
            O => \N__49240\,
            I => \N__48767\
        );

    \I__11620\ : SRMux
    port map (
            O => \N__49239\,
            I => \N__48767\
        );

    \I__11619\ : SRMux
    port map (
            O => \N__49238\,
            I => \N__48767\
        );

    \I__11618\ : SRMux
    port map (
            O => \N__49237\,
            I => \N__48767\
        );

    \I__11617\ : SRMux
    port map (
            O => \N__49236\,
            I => \N__48767\
        );

    \I__11616\ : SRMux
    port map (
            O => \N__49235\,
            I => \N__48767\
        );

    \I__11615\ : SRMux
    port map (
            O => \N__49234\,
            I => \N__48767\
        );

    \I__11614\ : SRMux
    port map (
            O => \N__49233\,
            I => \N__48767\
        );

    \I__11613\ : SRMux
    port map (
            O => \N__49232\,
            I => \N__48767\
        );

    \I__11612\ : SRMux
    port map (
            O => \N__49231\,
            I => \N__48767\
        );

    \I__11611\ : SRMux
    port map (
            O => \N__49230\,
            I => \N__48767\
        );

    \I__11610\ : SRMux
    port map (
            O => \N__49229\,
            I => \N__48767\
        );

    \I__11609\ : SRMux
    port map (
            O => \N__49228\,
            I => \N__48767\
        );

    \I__11608\ : SRMux
    port map (
            O => \N__49227\,
            I => \N__48767\
        );

    \I__11607\ : SRMux
    port map (
            O => \N__49226\,
            I => \N__48767\
        );

    \I__11606\ : SRMux
    port map (
            O => \N__49225\,
            I => \N__48767\
        );

    \I__11605\ : SRMux
    port map (
            O => \N__49224\,
            I => \N__48767\
        );

    \I__11604\ : SRMux
    port map (
            O => \N__49223\,
            I => \N__48767\
        );

    \I__11603\ : SRMux
    port map (
            O => \N__49222\,
            I => \N__48767\
        );

    \I__11602\ : SRMux
    port map (
            O => \N__49221\,
            I => \N__48767\
        );

    \I__11601\ : SRMux
    port map (
            O => \N__49220\,
            I => \N__48767\
        );

    \I__11600\ : SRMux
    port map (
            O => \N__49219\,
            I => \N__48767\
        );

    \I__11599\ : SRMux
    port map (
            O => \N__49218\,
            I => \N__48767\
        );

    \I__11598\ : SRMux
    port map (
            O => \N__49217\,
            I => \N__48767\
        );

    \I__11597\ : SRMux
    port map (
            O => \N__49216\,
            I => \N__48767\
        );

    \I__11596\ : SRMux
    port map (
            O => \N__49215\,
            I => \N__48767\
        );

    \I__11595\ : SRMux
    port map (
            O => \N__49214\,
            I => \N__48767\
        );

    \I__11594\ : SRMux
    port map (
            O => \N__49213\,
            I => \N__48767\
        );

    \I__11593\ : SRMux
    port map (
            O => \N__49212\,
            I => \N__48767\
        );

    \I__11592\ : SRMux
    port map (
            O => \N__49211\,
            I => \N__48767\
        );

    \I__11591\ : SRMux
    port map (
            O => \N__49210\,
            I => \N__48767\
        );

    \I__11590\ : SRMux
    port map (
            O => \N__49209\,
            I => \N__48767\
        );

    \I__11589\ : SRMux
    port map (
            O => \N__49208\,
            I => \N__48767\
        );

    \I__11588\ : SRMux
    port map (
            O => \N__49207\,
            I => \N__48767\
        );

    \I__11587\ : SRMux
    port map (
            O => \N__49206\,
            I => \N__48767\
        );

    \I__11586\ : SRMux
    port map (
            O => \N__49205\,
            I => \N__48767\
        );

    \I__11585\ : SRMux
    port map (
            O => \N__49204\,
            I => \N__48767\
        );

    \I__11584\ : SRMux
    port map (
            O => \N__49203\,
            I => \N__48767\
        );

    \I__11583\ : SRMux
    port map (
            O => \N__49202\,
            I => \N__48767\
        );

    \I__11582\ : SRMux
    port map (
            O => \N__49201\,
            I => \N__48767\
        );

    \I__11581\ : SRMux
    port map (
            O => \N__49200\,
            I => \N__48767\
        );

    \I__11580\ : SRMux
    port map (
            O => \N__49199\,
            I => \N__48767\
        );

    \I__11579\ : SRMux
    port map (
            O => \N__49198\,
            I => \N__48767\
        );

    \I__11578\ : SRMux
    port map (
            O => \N__49197\,
            I => \N__48767\
        );

    \I__11577\ : SRMux
    port map (
            O => \N__49196\,
            I => \N__48767\
        );

    \I__11576\ : SRMux
    port map (
            O => \N__49195\,
            I => \N__48767\
        );

    \I__11575\ : SRMux
    port map (
            O => \N__49194\,
            I => \N__48767\
        );

    \I__11574\ : SRMux
    port map (
            O => \N__49193\,
            I => \N__48767\
        );

    \I__11573\ : SRMux
    port map (
            O => \N__49192\,
            I => \N__48767\
        );

    \I__11572\ : SRMux
    port map (
            O => \N__49191\,
            I => \N__48767\
        );

    \I__11571\ : SRMux
    port map (
            O => \N__49190\,
            I => \N__48767\
        );

    \I__11570\ : SRMux
    port map (
            O => \N__49189\,
            I => \N__48767\
        );

    \I__11569\ : SRMux
    port map (
            O => \N__49188\,
            I => \N__48767\
        );

    \I__11568\ : SRMux
    port map (
            O => \N__49187\,
            I => \N__48767\
        );

    \I__11567\ : SRMux
    port map (
            O => \N__49186\,
            I => \N__48767\
        );

    \I__11566\ : SRMux
    port map (
            O => \N__49185\,
            I => \N__48767\
        );

    \I__11565\ : SRMux
    port map (
            O => \N__49184\,
            I => \N__48767\
        );

    \I__11564\ : SRMux
    port map (
            O => \N__49183\,
            I => \N__48767\
        );

    \I__11563\ : SRMux
    port map (
            O => \N__49182\,
            I => \N__48767\
        );

    \I__11562\ : SRMux
    port map (
            O => \N__49181\,
            I => \N__48767\
        );

    \I__11561\ : SRMux
    port map (
            O => \N__49180\,
            I => \N__48767\
        );

    \I__11560\ : SRMux
    port map (
            O => \N__49179\,
            I => \N__48767\
        );

    \I__11559\ : SRMux
    port map (
            O => \N__49178\,
            I => \N__48767\
        );

    \I__11558\ : SRMux
    port map (
            O => \N__49177\,
            I => \N__48767\
        );

    \I__11557\ : SRMux
    port map (
            O => \N__49176\,
            I => \N__48767\
        );

    \I__11556\ : SRMux
    port map (
            O => \N__49175\,
            I => \N__48767\
        );

    \I__11555\ : SRMux
    port map (
            O => \N__49174\,
            I => \N__48767\
        );

    \I__11554\ : SRMux
    port map (
            O => \N__49173\,
            I => \N__48767\
        );

    \I__11553\ : SRMux
    port map (
            O => \N__49172\,
            I => \N__48767\
        );

    \I__11552\ : SRMux
    port map (
            O => \N__49171\,
            I => \N__48767\
        );

    \I__11551\ : SRMux
    port map (
            O => \N__49170\,
            I => \N__48767\
        );

    \I__11550\ : SRMux
    port map (
            O => \N__49169\,
            I => \N__48767\
        );

    \I__11549\ : SRMux
    port map (
            O => \N__49168\,
            I => \N__48767\
        );

    \I__11548\ : SRMux
    port map (
            O => \N__49167\,
            I => \N__48767\
        );

    \I__11547\ : SRMux
    port map (
            O => \N__49166\,
            I => \N__48767\
        );

    \I__11546\ : SRMux
    port map (
            O => \N__49165\,
            I => \N__48767\
        );

    \I__11545\ : SRMux
    port map (
            O => \N__49164\,
            I => \N__48767\
        );

    \I__11544\ : SRMux
    port map (
            O => \N__49163\,
            I => \N__48767\
        );

    \I__11543\ : SRMux
    port map (
            O => \N__49162\,
            I => \N__48767\
        );

    \I__11542\ : SRMux
    port map (
            O => \N__49161\,
            I => \N__48767\
        );

    \I__11541\ : SRMux
    port map (
            O => \N__49160\,
            I => \N__48767\
        );

    \I__11540\ : SRMux
    port map (
            O => \N__49159\,
            I => \N__48767\
        );

    \I__11539\ : SRMux
    port map (
            O => \N__49158\,
            I => \N__48767\
        );

    \I__11538\ : SRMux
    port map (
            O => \N__49157\,
            I => \N__48767\
        );

    \I__11537\ : SRMux
    port map (
            O => \N__49156\,
            I => \N__48767\
        );

    \I__11536\ : SRMux
    port map (
            O => \N__49155\,
            I => \N__48767\
        );

    \I__11535\ : SRMux
    port map (
            O => \N__49154\,
            I => \N__48767\
        );

    \I__11534\ : SRMux
    port map (
            O => \N__49153\,
            I => \N__48767\
        );

    \I__11533\ : SRMux
    port map (
            O => \N__49152\,
            I => \N__48767\
        );

    \I__11532\ : SRMux
    port map (
            O => \N__49151\,
            I => \N__48767\
        );

    \I__11531\ : SRMux
    port map (
            O => \N__49150\,
            I => \N__48767\
        );

    \I__11530\ : SRMux
    port map (
            O => \N__49149\,
            I => \N__48767\
        );

    \I__11529\ : SRMux
    port map (
            O => \N__49148\,
            I => \N__48767\
        );

    \I__11528\ : SRMux
    port map (
            O => \N__49147\,
            I => \N__48767\
        );

    \I__11527\ : SRMux
    port map (
            O => \N__49146\,
            I => \N__48767\
        );

    \I__11526\ : SRMux
    port map (
            O => \N__49145\,
            I => \N__48767\
        );

    \I__11525\ : SRMux
    port map (
            O => \N__49144\,
            I => \N__48767\
        );

    \I__11524\ : SRMux
    port map (
            O => \N__49143\,
            I => \N__48767\
        );

    \I__11523\ : SRMux
    port map (
            O => \N__49142\,
            I => \N__48767\
        );

    \I__11522\ : SRMux
    port map (
            O => \N__49141\,
            I => \N__48767\
        );

    \I__11521\ : SRMux
    port map (
            O => \N__49140\,
            I => \N__48767\
        );

    \I__11520\ : SRMux
    port map (
            O => \N__49139\,
            I => \N__48767\
        );

    \I__11519\ : SRMux
    port map (
            O => \N__49138\,
            I => \N__48767\
        );

    \I__11518\ : SRMux
    port map (
            O => \N__49137\,
            I => \N__48767\
        );

    \I__11517\ : SRMux
    port map (
            O => \N__49136\,
            I => \N__48767\
        );

    \I__11516\ : SRMux
    port map (
            O => \N__49135\,
            I => \N__48767\
        );

    \I__11515\ : SRMux
    port map (
            O => \N__49134\,
            I => \N__48767\
        );

    \I__11514\ : SRMux
    port map (
            O => \N__49133\,
            I => \N__48767\
        );

    \I__11513\ : SRMux
    port map (
            O => \N__49132\,
            I => \N__48767\
        );

    \I__11512\ : SRMux
    port map (
            O => \N__49131\,
            I => \N__48767\
        );

    \I__11511\ : SRMux
    port map (
            O => \N__49130\,
            I => \N__48767\
        );

    \I__11510\ : SRMux
    port map (
            O => \N__49129\,
            I => \N__48767\
        );

    \I__11509\ : SRMux
    port map (
            O => \N__49128\,
            I => \N__48767\
        );

    \I__11508\ : SRMux
    port map (
            O => \N__49127\,
            I => \N__48767\
        );

    \I__11507\ : SRMux
    port map (
            O => \N__49126\,
            I => \N__48767\
        );

    \I__11506\ : SRMux
    port map (
            O => \N__49125\,
            I => \N__48767\
        );

    \I__11505\ : SRMux
    port map (
            O => \N__49124\,
            I => \N__48767\
        );

    \I__11504\ : SRMux
    port map (
            O => \N__49123\,
            I => \N__48767\
        );

    \I__11503\ : SRMux
    port map (
            O => \N__49122\,
            I => \N__48767\
        );

    \I__11502\ : SRMux
    port map (
            O => \N__49121\,
            I => \N__48767\
        );

    \I__11501\ : SRMux
    port map (
            O => \N__49120\,
            I => \N__48767\
        );

    \I__11500\ : SRMux
    port map (
            O => \N__49119\,
            I => \N__48767\
        );

    \I__11499\ : SRMux
    port map (
            O => \N__49118\,
            I => \N__48767\
        );

    \I__11498\ : SRMux
    port map (
            O => \N__49117\,
            I => \N__48767\
        );

    \I__11497\ : SRMux
    port map (
            O => \N__49116\,
            I => \N__48767\
        );

    \I__11496\ : SRMux
    port map (
            O => \N__49115\,
            I => \N__48767\
        );

    \I__11495\ : SRMux
    port map (
            O => \N__49114\,
            I => \N__48767\
        );

    \I__11494\ : SRMux
    port map (
            O => \N__49113\,
            I => \N__48767\
        );

    \I__11493\ : SRMux
    port map (
            O => \N__49112\,
            I => \N__48767\
        );

    \I__11492\ : SRMux
    port map (
            O => \N__49111\,
            I => \N__48767\
        );

    \I__11491\ : SRMux
    port map (
            O => \N__49110\,
            I => \N__48767\
        );

    \I__11490\ : SRMux
    port map (
            O => \N__49109\,
            I => \N__48767\
        );

    \I__11489\ : SRMux
    port map (
            O => \N__49108\,
            I => \N__48767\
        );

    \I__11488\ : SRMux
    port map (
            O => \N__49107\,
            I => \N__48767\
        );

    \I__11487\ : SRMux
    port map (
            O => \N__49106\,
            I => \N__48767\
        );

    \I__11486\ : SRMux
    port map (
            O => \N__49105\,
            I => \N__48767\
        );

    \I__11485\ : SRMux
    port map (
            O => \N__49104\,
            I => \N__48767\
        );

    \I__11484\ : SRMux
    port map (
            O => \N__49103\,
            I => \N__48767\
        );

    \I__11483\ : SRMux
    port map (
            O => \N__49102\,
            I => \N__48767\
        );

    \I__11482\ : SRMux
    port map (
            O => \N__49101\,
            I => \N__48767\
        );

    \I__11481\ : SRMux
    port map (
            O => \N__49100\,
            I => \N__48767\
        );

    \I__11480\ : SRMux
    port map (
            O => \N__49099\,
            I => \N__48767\
        );

    \I__11479\ : SRMux
    port map (
            O => \N__49098\,
            I => \N__48767\
        );

    \I__11478\ : SRMux
    port map (
            O => \N__49097\,
            I => \N__48767\
        );

    \I__11477\ : SRMux
    port map (
            O => \N__49096\,
            I => \N__48767\
        );

    \I__11476\ : SRMux
    port map (
            O => \N__49095\,
            I => \N__48767\
        );

    \I__11475\ : SRMux
    port map (
            O => \N__49094\,
            I => \N__48767\
        );

    \I__11474\ : SRMux
    port map (
            O => \N__49093\,
            I => \N__48767\
        );

    \I__11473\ : SRMux
    port map (
            O => \N__49092\,
            I => \N__48767\
        );

    \I__11472\ : SRMux
    port map (
            O => \N__49091\,
            I => \N__48767\
        );

    \I__11471\ : SRMux
    port map (
            O => \N__49090\,
            I => \N__48767\
        );

    \I__11470\ : SRMux
    port map (
            O => \N__49089\,
            I => \N__48767\
        );

    \I__11469\ : SRMux
    port map (
            O => \N__49088\,
            I => \N__48767\
        );

    \I__11468\ : GlobalMux
    port map (
            O => \N__48767\,
            I => \N__48764\
        );

    \I__11467\ : gio2CtrlBuf
    port map (
            O => \N__48764\,
            I => red_c_g
        );

    \I__11466\ : InMux
    port map (
            O => \N__48761\,
            I => \N__48754\
        );

    \I__11465\ : InMux
    port map (
            O => \N__48760\,
            I => \N__48754\
        );

    \I__11464\ : InMux
    port map (
            O => \N__48759\,
            I => \N__48751\
        );

    \I__11463\ : LocalMux
    port map (
            O => \N__48754\,
            I => \N__48748\
        );

    \I__11462\ : LocalMux
    port map (
            O => \N__48751\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__11461\ : Odrv12
    port map (
            O => \N__48748\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__11460\ : InMux
    port map (
            O => \N__48743\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__11459\ : CascadeMux
    port map (
            O => \N__48740\,
            I => \N__48736\
        );

    \I__11458\ : CascadeMux
    port map (
            O => \N__48739\,
            I => \N__48733\
        );

    \I__11457\ : InMux
    port map (
            O => \N__48736\,
            I => \N__48727\
        );

    \I__11456\ : InMux
    port map (
            O => \N__48733\,
            I => \N__48727\
        );

    \I__11455\ : InMux
    port map (
            O => \N__48732\,
            I => \N__48724\
        );

    \I__11454\ : LocalMux
    port map (
            O => \N__48727\,
            I => \N__48721\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__48724\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__11452\ : Odrv12
    port map (
            O => \N__48721\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__11451\ : InMux
    port map (
            O => \N__48716\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__11450\ : CascadeMux
    port map (
            O => \N__48713\,
            I => \N__48709\
        );

    \I__11449\ : InMux
    port map (
            O => \N__48712\,
            I => \N__48705\
        );

    \I__11448\ : InMux
    port map (
            O => \N__48709\,
            I => \N__48702\
        );

    \I__11447\ : InMux
    port map (
            O => \N__48708\,
            I => \N__48699\
        );

    \I__11446\ : LocalMux
    port map (
            O => \N__48705\,
            I => \N__48694\
        );

    \I__11445\ : LocalMux
    port map (
            O => \N__48702\,
            I => \N__48694\
        );

    \I__11444\ : LocalMux
    port map (
            O => \N__48699\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__11443\ : Odrv12
    port map (
            O => \N__48694\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__11442\ : InMux
    port map (
            O => \N__48689\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__11441\ : CascadeMux
    port map (
            O => \N__48686\,
            I => \N__48683\
        );

    \I__11440\ : InMux
    port map (
            O => \N__48683\,
            I => \N__48678\
        );

    \I__11439\ : InMux
    port map (
            O => \N__48682\,
            I => \N__48675\
        );

    \I__11438\ : InMux
    port map (
            O => \N__48681\,
            I => \N__48672\
        );

    \I__11437\ : LocalMux
    port map (
            O => \N__48678\,
            I => \N__48667\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__48675\,
            I => \N__48667\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__48672\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__11434\ : Odrv12
    port map (
            O => \N__48667\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__11433\ : InMux
    port map (
            O => \N__48662\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__11432\ : CascadeMux
    port map (
            O => \N__48659\,
            I => \N__48655\
        );

    \I__11431\ : CascadeMux
    port map (
            O => \N__48658\,
            I => \N__48652\
        );

    \I__11430\ : InMux
    port map (
            O => \N__48655\,
            I => \N__48647\
        );

    \I__11429\ : InMux
    port map (
            O => \N__48652\,
            I => \N__48647\
        );

    \I__11428\ : LocalMux
    port map (
            O => \N__48647\,
            I => \N__48643\
        );

    \I__11427\ : InMux
    port map (
            O => \N__48646\,
            I => \N__48640\
        );

    \I__11426\ : Span4Mux_v
    port map (
            O => \N__48643\,
            I => \N__48637\
        );

    \I__11425\ : LocalMux
    port map (
            O => \N__48640\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__11424\ : Odrv4
    port map (
            O => \N__48637\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__11423\ : InMux
    port map (
            O => \N__48632\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__11422\ : InMux
    port map (
            O => \N__48629\,
            I => \N__48622\
        );

    \I__11421\ : InMux
    port map (
            O => \N__48628\,
            I => \N__48622\
        );

    \I__11420\ : InMux
    port map (
            O => \N__48627\,
            I => \N__48619\
        );

    \I__11419\ : LocalMux
    port map (
            O => \N__48622\,
            I => \N__48616\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__48619\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__11417\ : Odrv12
    port map (
            O => \N__48616\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__11416\ : InMux
    port map (
            O => \N__48611\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__11415\ : CascadeMux
    port map (
            O => \N__48608\,
            I => \N__48605\
        );

    \I__11414\ : InMux
    port map (
            O => \N__48605\,
            I => \N__48601\
        );

    \I__11413\ : InMux
    port map (
            O => \N__48604\,
            I => \N__48598\
        );

    \I__11412\ : LocalMux
    port map (
            O => \N__48601\,
            I => \N__48592\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__48598\,
            I => \N__48592\
        );

    \I__11410\ : InMux
    port map (
            O => \N__48597\,
            I => \N__48589\
        );

    \I__11409\ : Span4Mux_v
    port map (
            O => \N__48592\,
            I => \N__48586\
        );

    \I__11408\ : LocalMux
    port map (
            O => \N__48589\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__11407\ : Odrv4
    port map (
            O => \N__48586\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__11406\ : InMux
    port map (
            O => \N__48581\,
            I => \bfn_18_26_0_\
        );

    \I__11405\ : CascadeMux
    port map (
            O => \N__48578\,
            I => \N__48574\
        );

    \I__11404\ : InMux
    port map (
            O => \N__48577\,
            I => \N__48571\
        );

    \I__11403\ : InMux
    port map (
            O => \N__48574\,
            I => \N__48568\
        );

    \I__11402\ : LocalMux
    port map (
            O => \N__48571\,
            I => \N__48562\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__48568\,
            I => \N__48562\
        );

    \I__11400\ : InMux
    port map (
            O => \N__48567\,
            I => \N__48559\
        );

    \I__11399\ : Span4Mux_v
    port map (
            O => \N__48562\,
            I => \N__48556\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__48559\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__11397\ : Odrv4
    port map (
            O => \N__48556\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__11396\ : InMux
    port map (
            O => \N__48551\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__11395\ : CascadeMux
    port map (
            O => \N__48548\,
            I => \N__48545\
        );

    \I__11394\ : InMux
    port map (
            O => \N__48545\,
            I => \N__48541\
        );

    \I__11393\ : InMux
    port map (
            O => \N__48544\,
            I => \N__48538\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__48541\,
            I => \N__48532\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__48538\,
            I => \N__48532\
        );

    \I__11390\ : InMux
    port map (
            O => \N__48537\,
            I => \N__48529\
        );

    \I__11389\ : Span4Mux_v
    port map (
            O => \N__48532\,
            I => \N__48526\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__48529\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__11387\ : Odrv4
    port map (
            O => \N__48526\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__11386\ : InMux
    port map (
            O => \N__48521\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__11385\ : InMux
    port map (
            O => \N__48518\,
            I => \N__48512\
        );

    \I__11384\ : InMux
    port map (
            O => \N__48517\,
            I => \N__48512\
        );

    \I__11383\ : LocalMux
    port map (
            O => \N__48512\,
            I => \N__48508\
        );

    \I__11382\ : InMux
    port map (
            O => \N__48511\,
            I => \N__48505\
        );

    \I__11381\ : Span4Mux_h
    port map (
            O => \N__48508\,
            I => \N__48502\
        );

    \I__11380\ : LocalMux
    port map (
            O => \N__48505\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__11379\ : Odrv4
    port map (
            O => \N__48502\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__11378\ : InMux
    port map (
            O => \N__48497\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__11377\ : InMux
    port map (
            O => \N__48494\,
            I => \N__48488\
        );

    \I__11376\ : InMux
    port map (
            O => \N__48493\,
            I => \N__48488\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__48488\,
            I => \N__48484\
        );

    \I__11374\ : InMux
    port map (
            O => \N__48487\,
            I => \N__48481\
        );

    \I__11373\ : Span4Mux_h
    port map (
            O => \N__48484\,
            I => \N__48478\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__48481\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__11371\ : Odrv4
    port map (
            O => \N__48478\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__11370\ : InMux
    port map (
            O => \N__48473\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__11369\ : CascadeMux
    port map (
            O => \N__48470\,
            I => \N__48466\
        );

    \I__11368\ : CascadeMux
    port map (
            O => \N__48469\,
            I => \N__48463\
        );

    \I__11367\ : InMux
    port map (
            O => \N__48466\,
            I => \N__48458\
        );

    \I__11366\ : InMux
    port map (
            O => \N__48463\,
            I => \N__48458\
        );

    \I__11365\ : LocalMux
    port map (
            O => \N__48458\,
            I => \N__48454\
        );

    \I__11364\ : InMux
    port map (
            O => \N__48457\,
            I => \N__48451\
        );

    \I__11363\ : Span4Mux_v
    port map (
            O => \N__48454\,
            I => \N__48448\
        );

    \I__11362\ : LocalMux
    port map (
            O => \N__48451\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__11361\ : Odrv4
    port map (
            O => \N__48448\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__11360\ : InMux
    port map (
            O => \N__48443\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__11359\ : CascadeMux
    port map (
            O => \N__48440\,
            I => \N__48436\
        );

    \I__11358\ : CascadeMux
    port map (
            O => \N__48439\,
            I => \N__48433\
        );

    \I__11357\ : InMux
    port map (
            O => \N__48436\,
            I => \N__48428\
        );

    \I__11356\ : InMux
    port map (
            O => \N__48433\,
            I => \N__48428\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__48428\,
            I => \N__48424\
        );

    \I__11354\ : InMux
    port map (
            O => \N__48427\,
            I => \N__48421\
        );

    \I__11353\ : Span4Mux_h
    port map (
            O => \N__48424\,
            I => \N__48418\
        );

    \I__11352\ : LocalMux
    port map (
            O => \N__48421\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__11351\ : Odrv4
    port map (
            O => \N__48418\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__11350\ : InMux
    port map (
            O => \N__48413\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__11349\ : InMux
    port map (
            O => \N__48410\,
            I => \N__48404\
        );

    \I__11348\ : InMux
    port map (
            O => \N__48409\,
            I => \N__48404\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__48404\,
            I => \N__48400\
        );

    \I__11346\ : InMux
    port map (
            O => \N__48403\,
            I => \N__48397\
        );

    \I__11345\ : Span4Mux_v
    port map (
            O => \N__48400\,
            I => \N__48394\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__48397\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__11343\ : Odrv4
    port map (
            O => \N__48394\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__11342\ : InMux
    port map (
            O => \N__48389\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__11341\ : CascadeMux
    port map (
            O => \N__48386\,
            I => \N__48383\
        );

    \I__11340\ : InMux
    port map (
            O => \N__48383\,
            I => \N__48379\
        );

    \I__11339\ : InMux
    port map (
            O => \N__48382\,
            I => \N__48376\
        );

    \I__11338\ : LocalMux
    port map (
            O => \N__48379\,
            I => \N__48370\
        );

    \I__11337\ : LocalMux
    port map (
            O => \N__48376\,
            I => \N__48370\
        );

    \I__11336\ : InMux
    port map (
            O => \N__48375\,
            I => \N__48367\
        );

    \I__11335\ : Span4Mux_v
    port map (
            O => \N__48370\,
            I => \N__48364\
        );

    \I__11334\ : LocalMux
    port map (
            O => \N__48367\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__11333\ : Odrv4
    port map (
            O => \N__48364\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__11332\ : InMux
    port map (
            O => \N__48359\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__11331\ : CascadeMux
    port map (
            O => \N__48356\,
            I => \N__48352\
        );

    \I__11330\ : CascadeMux
    port map (
            O => \N__48355\,
            I => \N__48349\
        );

    \I__11329\ : InMux
    port map (
            O => \N__48352\,
            I => \N__48346\
        );

    \I__11328\ : InMux
    port map (
            O => \N__48349\,
            I => \N__48343\
        );

    \I__11327\ : LocalMux
    port map (
            O => \N__48346\,
            I => \N__48337\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__48343\,
            I => \N__48337\
        );

    \I__11325\ : InMux
    port map (
            O => \N__48342\,
            I => \N__48334\
        );

    \I__11324\ : Span4Mux_v
    port map (
            O => \N__48337\,
            I => \N__48331\
        );

    \I__11323\ : LocalMux
    port map (
            O => \N__48334\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__11322\ : Odrv4
    port map (
            O => \N__48331\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__11321\ : InMux
    port map (
            O => \N__48326\,
            I => \bfn_18_25_0_\
        );

    \I__11320\ : InMux
    port map (
            O => \N__48323\,
            I => \N__48319\
        );

    \I__11319\ : InMux
    port map (
            O => \N__48322\,
            I => \N__48316\
        );

    \I__11318\ : LocalMux
    port map (
            O => \N__48319\,
            I => \N__48310\
        );

    \I__11317\ : LocalMux
    port map (
            O => \N__48316\,
            I => \N__48310\
        );

    \I__11316\ : InMux
    port map (
            O => \N__48315\,
            I => \N__48307\
        );

    \I__11315\ : Span4Mux_v
    port map (
            O => \N__48310\,
            I => \N__48304\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__48307\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__11313\ : Odrv4
    port map (
            O => \N__48304\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__11312\ : InMux
    port map (
            O => \N__48299\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__11311\ : InMux
    port map (
            O => \N__48296\,
            I => \N__48293\
        );

    \I__11310\ : LocalMux
    port map (
            O => \N__48293\,
            I => \N__48289\
        );

    \I__11309\ : CascadeMux
    port map (
            O => \N__48292\,
            I => \N__48286\
        );

    \I__11308\ : Span4Mux_v
    port map (
            O => \N__48289\,
            I => \N__48283\
        );

    \I__11307\ : InMux
    port map (
            O => \N__48286\,
            I => \N__48280\
        );

    \I__11306\ : Span4Mux_v
    port map (
            O => \N__48283\,
            I => \N__48277\
        );

    \I__11305\ : LocalMux
    port map (
            O => \N__48280\,
            I => \N__48273\
        );

    \I__11304\ : Span4Mux_v
    port map (
            O => \N__48277\,
            I => \N__48270\
        );

    \I__11303\ : InMux
    port map (
            O => \N__48276\,
            I => \N__48267\
        );

    \I__11302\ : Span4Mux_h
    port map (
            O => \N__48273\,
            I => \N__48264\
        );

    \I__11301\ : Odrv4
    port map (
            O => \N__48270\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__48267\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__11299\ : Odrv4
    port map (
            O => \N__48264\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__11298\ : InMux
    port map (
            O => \N__48257\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__11297\ : InMux
    port map (
            O => \N__48254\,
            I => \N__48247\
        );

    \I__11296\ : InMux
    port map (
            O => \N__48253\,
            I => \N__48247\
        );

    \I__11295\ : InMux
    port map (
            O => \N__48252\,
            I => \N__48244\
        );

    \I__11294\ : LocalMux
    port map (
            O => \N__48247\,
            I => \N__48241\
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__48244\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__11292\ : Odrv12
    port map (
            O => \N__48241\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__11291\ : InMux
    port map (
            O => \N__48236\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__11290\ : InMux
    port map (
            O => \N__48233\,
            I => \N__48226\
        );

    \I__11289\ : InMux
    port map (
            O => \N__48232\,
            I => \N__48226\
        );

    \I__11288\ : InMux
    port map (
            O => \N__48231\,
            I => \N__48223\
        );

    \I__11287\ : LocalMux
    port map (
            O => \N__48226\,
            I => \N__48220\
        );

    \I__11286\ : LocalMux
    port map (
            O => \N__48223\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__11285\ : Odrv12
    port map (
            O => \N__48220\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__11284\ : InMux
    port map (
            O => \N__48215\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__11283\ : CascadeMux
    port map (
            O => \N__48212\,
            I => \N__48208\
        );

    \I__11282\ : InMux
    port map (
            O => \N__48211\,
            I => \N__48205\
        );

    \I__11281\ : InMux
    port map (
            O => \N__48208\,
            I => \N__48202\
        );

    \I__11280\ : LocalMux
    port map (
            O => \N__48205\,
            I => \N__48196\
        );

    \I__11279\ : LocalMux
    port map (
            O => \N__48202\,
            I => \N__48196\
        );

    \I__11278\ : InMux
    port map (
            O => \N__48201\,
            I => \N__48193\
        );

    \I__11277\ : Span4Mux_h
    port map (
            O => \N__48196\,
            I => \N__48190\
        );

    \I__11276\ : LocalMux
    port map (
            O => \N__48193\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__11275\ : Odrv4
    port map (
            O => \N__48190\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__11274\ : InMux
    port map (
            O => \N__48185\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__11273\ : CascadeMux
    port map (
            O => \N__48182\,
            I => \N__48178\
        );

    \I__11272\ : InMux
    port map (
            O => \N__48181\,
            I => \N__48175\
        );

    \I__11271\ : InMux
    port map (
            O => \N__48178\,
            I => \N__48172\
        );

    \I__11270\ : LocalMux
    port map (
            O => \N__48175\,
            I => \N__48166\
        );

    \I__11269\ : LocalMux
    port map (
            O => \N__48172\,
            I => \N__48166\
        );

    \I__11268\ : InMux
    port map (
            O => \N__48171\,
            I => \N__48163\
        );

    \I__11267\ : Span4Mux_h
    port map (
            O => \N__48166\,
            I => \N__48160\
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__48163\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__11265\ : Odrv4
    port map (
            O => \N__48160\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__11264\ : InMux
    port map (
            O => \N__48155\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__11263\ : CascadeMux
    port map (
            O => \N__48152\,
            I => \N__48148\
        );

    \I__11262\ : CascadeMux
    port map (
            O => \N__48151\,
            I => \N__48145\
        );

    \I__11261\ : InMux
    port map (
            O => \N__48148\,
            I => \N__48140\
        );

    \I__11260\ : InMux
    port map (
            O => \N__48145\,
            I => \N__48140\
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__48140\,
            I => \N__48136\
        );

    \I__11258\ : InMux
    port map (
            O => \N__48139\,
            I => \N__48133\
        );

    \I__11257\ : Span4Mux_v
    port map (
            O => \N__48136\,
            I => \N__48130\
        );

    \I__11256\ : LocalMux
    port map (
            O => \N__48133\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__11255\ : Odrv4
    port map (
            O => \N__48130\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__11254\ : InMux
    port map (
            O => \N__48125\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__11253\ : CascadeMux
    port map (
            O => \N__48122\,
            I => \N__48118\
        );

    \I__11252\ : CascadeMux
    port map (
            O => \N__48121\,
            I => \N__48115\
        );

    \I__11251\ : InMux
    port map (
            O => \N__48118\,
            I => \N__48110\
        );

    \I__11250\ : InMux
    port map (
            O => \N__48115\,
            I => \N__48110\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__48110\,
            I => \N__48106\
        );

    \I__11248\ : InMux
    port map (
            O => \N__48109\,
            I => \N__48103\
        );

    \I__11247\ : Span4Mux_v
    port map (
            O => \N__48106\,
            I => \N__48100\
        );

    \I__11246\ : LocalMux
    port map (
            O => \N__48103\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__11245\ : Odrv4
    port map (
            O => \N__48100\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__11244\ : InMux
    port map (
            O => \N__48095\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__11243\ : CascadeMux
    port map (
            O => \N__48092\,
            I => \N__48089\
        );

    \I__11242\ : InMux
    port map (
            O => \N__48089\,
            I => \N__48085\
        );

    \I__11241\ : InMux
    port map (
            O => \N__48088\,
            I => \N__48082\
        );

    \I__11240\ : LocalMux
    port map (
            O => \N__48085\,
            I => \N__48076\
        );

    \I__11239\ : LocalMux
    port map (
            O => \N__48082\,
            I => \N__48076\
        );

    \I__11238\ : InMux
    port map (
            O => \N__48081\,
            I => \N__48073\
        );

    \I__11237\ : Span4Mux_v
    port map (
            O => \N__48076\,
            I => \N__48070\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__48073\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__11235\ : Odrv4
    port map (
            O => \N__48070\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__11234\ : InMux
    port map (
            O => \N__48065\,
            I => \bfn_18_24_0_\
        );

    \I__11233\ : InMux
    port map (
            O => \N__48062\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__11232\ : CascadeMux
    port map (
            O => \N__48059\,
            I => \N__48056\
        );

    \I__11231\ : InMux
    port map (
            O => \N__48056\,
            I => \N__48052\
        );

    \I__11230\ : CascadeMux
    port map (
            O => \N__48055\,
            I => \N__48049\
        );

    \I__11229\ : LocalMux
    port map (
            O => \N__48052\,
            I => \N__48046\
        );

    \I__11228\ : InMux
    port map (
            O => \N__48049\,
            I => \N__48043\
        );

    \I__11227\ : Span4Mux_h
    port map (
            O => \N__48046\,
            I => \N__48037\
        );

    \I__11226\ : LocalMux
    port map (
            O => \N__48043\,
            I => \N__48037\
        );

    \I__11225\ : InMux
    port map (
            O => \N__48042\,
            I => \N__48034\
        );

    \I__11224\ : Span4Mux_h
    port map (
            O => \N__48037\,
            I => \N__48030\
        );

    \I__11223\ : LocalMux
    port map (
            O => \N__48034\,
            I => \N__48027\
        );

    \I__11222\ : InMux
    port map (
            O => \N__48033\,
            I => \N__48024\
        );

    \I__11221\ : Odrv4
    port map (
            O => \N__48030\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__11220\ : Odrv4
    port map (
            O => \N__48027\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__11219\ : LocalMux
    port map (
            O => \N__48024\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__11218\ : InMux
    port map (
            O => \N__48017\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__11217\ : CascadeMux
    port map (
            O => \N__48014\,
            I => \N__48011\
        );

    \I__11216\ : InMux
    port map (
            O => \N__48011\,
            I => \N__48007\
        );

    \I__11215\ : InMux
    port map (
            O => \N__48010\,
            I => \N__48004\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__48007\,
            I => \N__48000\
        );

    \I__11213\ : LocalMux
    port map (
            O => \N__48004\,
            I => \N__47997\
        );

    \I__11212\ : InMux
    port map (
            O => \N__48003\,
            I => \N__47994\
        );

    \I__11211\ : Span4Mux_h
    port map (
            O => \N__48000\,
            I => \N__47990\
        );

    \I__11210\ : Span4Mux_h
    port map (
            O => \N__47997\,
            I => \N__47987\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__47994\,
            I => \N__47984\
        );

    \I__11208\ : InMux
    port map (
            O => \N__47993\,
            I => \N__47981\
        );

    \I__11207\ : Odrv4
    port map (
            O => \N__47990\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__11206\ : Odrv4
    port map (
            O => \N__47987\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__11205\ : Odrv4
    port map (
            O => \N__47984\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__11204\ : LocalMux
    port map (
            O => \N__47981\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__11203\ : InMux
    port map (
            O => \N__47972\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__11202\ : CascadeMux
    port map (
            O => \N__47969\,
            I => \N__47965\
        );

    \I__11201\ : InMux
    port map (
            O => \N__47968\,
            I => \N__47962\
        );

    \I__11200\ : InMux
    port map (
            O => \N__47965\,
            I => \N__47959\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__47962\,
            I => \N__47956\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__47959\,
            I => \N__47952\
        );

    \I__11197\ : Span4Mux_h
    port map (
            O => \N__47956\,
            I => \N__47949\
        );

    \I__11196\ : InMux
    port map (
            O => \N__47955\,
            I => \N__47946\
        );

    \I__11195\ : Span4Mux_h
    port map (
            O => \N__47952\,
            I => \N__47942\
        );

    \I__11194\ : Span4Mux_v
    port map (
            O => \N__47949\,
            I => \N__47937\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__47946\,
            I => \N__47937\
        );

    \I__11192\ : InMux
    port map (
            O => \N__47945\,
            I => \N__47934\
        );

    \I__11191\ : Odrv4
    port map (
            O => \N__47942\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__11190\ : Odrv4
    port map (
            O => \N__47937\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__47934\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__11188\ : InMux
    port map (
            O => \N__47927\,
            I => \bfn_18_22_0_\
        );

    \I__11187\ : CascadeMux
    port map (
            O => \N__47924\,
            I => \N__47920\
        );

    \I__11186\ : CascadeMux
    port map (
            O => \N__47923\,
            I => \N__47917\
        );

    \I__11185\ : InMux
    port map (
            O => \N__47920\,
            I => \N__47914\
        );

    \I__11184\ : InMux
    port map (
            O => \N__47917\,
            I => \N__47911\
        );

    \I__11183\ : LocalMux
    port map (
            O => \N__47914\,
            I => \N__47907\
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__47911\,
            I => \N__47904\
        );

    \I__11181\ : InMux
    port map (
            O => \N__47910\,
            I => \N__47901\
        );

    \I__11180\ : Span4Mux_h
    port map (
            O => \N__47907\,
            I => \N__47897\
        );

    \I__11179\ : Span4Mux_h
    port map (
            O => \N__47904\,
            I => \N__47894\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__47901\,
            I => \N__47891\
        );

    \I__11177\ : InMux
    port map (
            O => \N__47900\,
            I => \N__47888\
        );

    \I__11176\ : Odrv4
    port map (
            O => \N__47897\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11175\ : Odrv4
    port map (
            O => \N__47894\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11174\ : Odrv4
    port map (
            O => \N__47891\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11173\ : LocalMux
    port map (
            O => \N__47888\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11172\ : InMux
    port map (
            O => \N__47879\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__11171\ : InMux
    port map (
            O => \N__47876\,
            I => \N__47872\
        );

    \I__11170\ : InMux
    port map (
            O => \N__47875\,
            I => \N__47869\
        );

    \I__11169\ : LocalMux
    port map (
            O => \N__47872\,
            I => \N__47863\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__47869\,
            I => \N__47863\
        );

    \I__11167\ : InMux
    port map (
            O => \N__47868\,
            I => \N__47860\
        );

    \I__11166\ : Span4Mux_v
    port map (
            O => \N__47863\,
            I => \N__47856\
        );

    \I__11165\ : LocalMux
    port map (
            O => \N__47860\,
            I => \N__47853\
        );

    \I__11164\ : InMux
    port map (
            O => \N__47859\,
            I => \N__47850\
        );

    \I__11163\ : Odrv4
    port map (
            O => \N__47856\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__11162\ : Odrv4
    port map (
            O => \N__47853\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__11161\ : LocalMux
    port map (
            O => \N__47850\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__11160\ : InMux
    port map (
            O => \N__47843\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__11159\ : CascadeMux
    port map (
            O => \N__47840\,
            I => \N__47837\
        );

    \I__11158\ : InMux
    port map (
            O => \N__47837\,
            I => \N__47833\
        );

    \I__11157\ : CascadeMux
    port map (
            O => \N__47836\,
            I => \N__47830\
        );

    \I__11156\ : LocalMux
    port map (
            O => \N__47833\,
            I => \N__47827\
        );

    \I__11155\ : InMux
    port map (
            O => \N__47830\,
            I => \N__47824\
        );

    \I__11154\ : Span4Mux_v
    port map (
            O => \N__47827\,
            I => \N__47818\
        );

    \I__11153\ : LocalMux
    port map (
            O => \N__47824\,
            I => \N__47818\
        );

    \I__11152\ : InMux
    port map (
            O => \N__47823\,
            I => \N__47815\
        );

    \I__11151\ : Span4Mux_h
    port map (
            O => \N__47818\,
            I => \N__47811\
        );

    \I__11150\ : LocalMux
    port map (
            O => \N__47815\,
            I => \N__47808\
        );

    \I__11149\ : InMux
    port map (
            O => \N__47814\,
            I => \N__47805\
        );

    \I__11148\ : Odrv4
    port map (
            O => \N__47811\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__11147\ : Odrv4
    port map (
            O => \N__47808\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__11146\ : LocalMux
    port map (
            O => \N__47805\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__11145\ : InMux
    port map (
            O => \N__47798\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__11144\ : CEMux
    port map (
            O => \N__47795\,
            I => \N__47771\
        );

    \I__11143\ : CEMux
    port map (
            O => \N__47794\,
            I => \N__47771\
        );

    \I__11142\ : CEMux
    port map (
            O => \N__47793\,
            I => \N__47771\
        );

    \I__11141\ : CEMux
    port map (
            O => \N__47792\,
            I => \N__47771\
        );

    \I__11140\ : CEMux
    port map (
            O => \N__47791\,
            I => \N__47771\
        );

    \I__11139\ : CEMux
    port map (
            O => \N__47790\,
            I => \N__47771\
        );

    \I__11138\ : CEMux
    port map (
            O => \N__47789\,
            I => \N__47771\
        );

    \I__11137\ : CEMux
    port map (
            O => \N__47788\,
            I => \N__47771\
        );

    \I__11136\ : GlobalMux
    port map (
            O => \N__47771\,
            I => \N__47768\
        );

    \I__11135\ : gio2CtrlBuf
    port map (
            O => \N__47768\,
            I => \current_shift_inst.timer_s1.N_161_i_g\
        );

    \I__11134\ : InMux
    port map (
            O => \N__47765\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__11133\ : InMux
    port map (
            O => \N__47762\,
            I => \N__47759\
        );

    \I__11132\ : LocalMux
    port map (
            O => \N__47759\,
            I => \N__47754\
        );

    \I__11131\ : InMux
    port map (
            O => \N__47758\,
            I => \N__47751\
        );

    \I__11130\ : InMux
    port map (
            O => \N__47757\,
            I => \N__47748\
        );

    \I__11129\ : Span4Mux_v
    port map (
            O => \N__47754\,
            I => \N__47745\
        );

    \I__11128\ : LocalMux
    port map (
            O => \N__47751\,
            I => \N__47742\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__47748\,
            I => \N__47739\
        );

    \I__11126\ : Span4Mux_v
    port map (
            O => \N__47745\,
            I => \N__47736\
        );

    \I__11125\ : Span12Mux_h
    port map (
            O => \N__47742\,
            I => \N__47731\
        );

    \I__11124\ : Span12Mux_v
    port map (
            O => \N__47739\,
            I => \N__47731\
        );

    \I__11123\ : Odrv4
    port map (
            O => \N__47736\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__11122\ : Odrv12
    port map (
            O => \N__47731\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__11121\ : InMux
    port map (
            O => \N__47726\,
            I => \N__47723\
        );

    \I__11120\ : LocalMux
    port map (
            O => \N__47723\,
            I => \N__47719\
        );

    \I__11119\ : CascadeMux
    port map (
            O => \N__47722\,
            I => \N__47716\
        );

    \I__11118\ : Span4Mux_h
    port map (
            O => \N__47719\,
            I => \N__47713\
        );

    \I__11117\ : InMux
    port map (
            O => \N__47716\,
            I => \N__47709\
        );

    \I__11116\ : Span4Mux_v
    port map (
            O => \N__47713\,
            I => \N__47706\
        );

    \I__11115\ : InMux
    port map (
            O => \N__47712\,
            I => \N__47703\
        );

    \I__11114\ : LocalMux
    port map (
            O => \N__47709\,
            I => \N__47700\
        );

    \I__11113\ : Odrv4
    port map (
            O => \N__47706\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__47703\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__11111\ : Odrv12
    port map (
            O => \N__47700\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__11110\ : InMux
    port map (
            O => \N__47693\,
            I => \bfn_18_23_0_\
        );

    \I__11109\ : CascadeMux
    port map (
            O => \N__47690\,
            I => \N__47686\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47689\,
            I => \N__47682\
        );

    \I__11107\ : InMux
    port map (
            O => \N__47686\,
            I => \N__47679\
        );

    \I__11106\ : InMux
    port map (
            O => \N__47685\,
            I => \N__47676\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__47682\,
            I => \N__47672\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__47679\,
            I => \N__47667\
        );

    \I__11103\ : LocalMux
    port map (
            O => \N__47676\,
            I => \N__47667\
        );

    \I__11102\ : InMux
    port map (
            O => \N__47675\,
            I => \N__47664\
        );

    \I__11101\ : Span12Mux_h
    port map (
            O => \N__47672\,
            I => \N__47661\
        );

    \I__11100\ : Span4Mux_v
    port map (
            O => \N__47667\,
            I => \N__47656\
        );

    \I__11099\ : LocalMux
    port map (
            O => \N__47664\,
            I => \N__47656\
        );

    \I__11098\ : Odrv12
    port map (
            O => \N__47661\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__11097\ : Odrv4
    port map (
            O => \N__47656\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__11096\ : InMux
    port map (
            O => \N__47651\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__11095\ : CascadeMux
    port map (
            O => \N__47648\,
            I => \N__47645\
        );

    \I__11094\ : InMux
    port map (
            O => \N__47645\,
            I => \N__47640\
        );

    \I__11093\ : InMux
    port map (
            O => \N__47644\,
            I => \N__47637\
        );

    \I__11092\ : InMux
    port map (
            O => \N__47643\,
            I => \N__47634\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__47640\,
            I => \N__47631\
        );

    \I__11090\ : LocalMux
    port map (
            O => \N__47637\,
            I => \N__47628\
        );

    \I__11089\ : LocalMux
    port map (
            O => \N__47634\,
            I => \N__47625\
        );

    \I__11088\ : Sp12to4
    port map (
            O => \N__47631\,
            I => \N__47621\
        );

    \I__11087\ : Span4Mux_v
    port map (
            O => \N__47628\,
            I => \N__47618\
        );

    \I__11086\ : Span4Mux_v
    port map (
            O => \N__47625\,
            I => \N__47615\
        );

    \I__11085\ : InMux
    port map (
            O => \N__47624\,
            I => \N__47612\
        );

    \I__11084\ : Odrv12
    port map (
            O => \N__47621\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__11083\ : Odrv4
    port map (
            O => \N__47618\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__11082\ : Odrv4
    port map (
            O => \N__47615\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__47612\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__11080\ : InMux
    port map (
            O => \N__47603\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__11079\ : CascadeMux
    port map (
            O => \N__47600\,
            I => \N__47596\
        );

    \I__11078\ : InMux
    port map (
            O => \N__47599\,
            I => \N__47592\
        );

    \I__11077\ : InMux
    port map (
            O => \N__47596\,
            I => \N__47589\
        );

    \I__11076\ : InMux
    port map (
            O => \N__47595\,
            I => \N__47586\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__47592\,
            I => \N__47581\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__47589\,
            I => \N__47581\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__47586\,
            I => \N__47578\
        );

    \I__11072\ : Span4Mux_h
    port map (
            O => \N__47581\,
            I => \N__47574\
        );

    \I__11071\ : Span4Mux_h
    port map (
            O => \N__47578\,
            I => \N__47571\
        );

    \I__11070\ : InMux
    port map (
            O => \N__47577\,
            I => \N__47568\
        );

    \I__11069\ : Odrv4
    port map (
            O => \N__47574\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__11068\ : Odrv4
    port map (
            O => \N__47571\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__11067\ : LocalMux
    port map (
            O => \N__47568\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__11066\ : InMux
    port map (
            O => \N__47561\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__11065\ : CascadeMux
    port map (
            O => \N__47558\,
            I => \N__47555\
        );

    \I__11064\ : InMux
    port map (
            O => \N__47555\,
            I => \N__47551\
        );

    \I__11063\ : InMux
    port map (
            O => \N__47554\,
            I => \N__47548\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__47551\,
            I => \N__47545\
        );

    \I__11061\ : LocalMux
    port map (
            O => \N__47548\,
            I => \N__47542\
        );

    \I__11060\ : Span4Mux_v
    port map (
            O => \N__47545\,
            I => \N__47537\
        );

    \I__11059\ : Span12Mux_v
    port map (
            O => \N__47542\,
            I => \N__47534\
        );

    \I__11058\ : InMux
    port map (
            O => \N__47541\,
            I => \N__47531\
        );

    \I__11057\ : InMux
    port map (
            O => \N__47540\,
            I => \N__47528\
        );

    \I__11056\ : Odrv4
    port map (
            O => \N__47537\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__11055\ : Odrv12
    port map (
            O => \N__47534\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__47531\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__11053\ : LocalMux
    port map (
            O => \N__47528\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__11052\ : InMux
    port map (
            O => \N__47519\,
            I => \bfn_18_21_0_\
        );

    \I__11051\ : CascadeMux
    port map (
            O => \N__47516\,
            I => \N__47513\
        );

    \I__11050\ : InMux
    port map (
            O => \N__47513\,
            I => \N__47509\
        );

    \I__11049\ : CascadeMux
    port map (
            O => \N__47512\,
            I => \N__47506\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__47509\,
            I => \N__47503\
        );

    \I__11047\ : InMux
    port map (
            O => \N__47506\,
            I => \N__47500\
        );

    \I__11046\ : Span4Mux_h
    port map (
            O => \N__47503\,
            I => \N__47495\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__47500\,
            I => \N__47495\
        );

    \I__11044\ : Span4Mux_v
    port map (
            O => \N__47495\,
            I => \N__47490\
        );

    \I__11043\ : InMux
    port map (
            O => \N__47494\,
            I => \N__47487\
        );

    \I__11042\ : InMux
    port map (
            O => \N__47493\,
            I => \N__47484\
        );

    \I__11041\ : Odrv4
    port map (
            O => \N__47490\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__47487\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__47484\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__11038\ : InMux
    port map (
            O => \N__47477\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__11037\ : CascadeMux
    port map (
            O => \N__47474\,
            I => \N__47470\
        );

    \I__11036\ : CascadeMux
    port map (
            O => \N__47473\,
            I => \N__47467\
        );

    \I__11035\ : InMux
    port map (
            O => \N__47470\,
            I => \N__47464\
        );

    \I__11034\ : InMux
    port map (
            O => \N__47467\,
            I => \N__47461\
        );

    \I__11033\ : LocalMux
    port map (
            O => \N__47464\,
            I => \N__47455\
        );

    \I__11032\ : LocalMux
    port map (
            O => \N__47461\,
            I => \N__47455\
        );

    \I__11031\ : InMux
    port map (
            O => \N__47460\,
            I => \N__47452\
        );

    \I__11030\ : Span4Mux_v
    port map (
            O => \N__47455\,
            I => \N__47447\
        );

    \I__11029\ : LocalMux
    port map (
            O => \N__47452\,
            I => \N__47447\
        );

    \I__11028\ : Span4Mux_h
    port map (
            O => \N__47447\,
            I => \N__47443\
        );

    \I__11027\ : InMux
    port map (
            O => \N__47446\,
            I => \N__47440\
        );

    \I__11026\ : Odrv4
    port map (
            O => \N__47443\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__47440\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__11024\ : InMux
    port map (
            O => \N__47435\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__11023\ : CascadeMux
    port map (
            O => \N__47432\,
            I => \N__47428\
        );

    \I__11022\ : InMux
    port map (
            O => \N__47431\,
            I => \N__47425\
        );

    \I__11021\ : InMux
    port map (
            O => \N__47428\,
            I => \N__47422\
        );

    \I__11020\ : LocalMux
    port map (
            O => \N__47425\,
            I => \N__47418\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__47422\,
            I => \N__47415\
        );

    \I__11018\ : InMux
    port map (
            O => \N__47421\,
            I => \N__47412\
        );

    \I__11017\ : Span4Mux_h
    port map (
            O => \N__47418\,
            I => \N__47409\
        );

    \I__11016\ : Span4Mux_h
    port map (
            O => \N__47415\,
            I => \N__47405\
        );

    \I__11015\ : LocalMux
    port map (
            O => \N__47412\,
            I => \N__47402\
        );

    \I__11014\ : Span4Mux_v
    port map (
            O => \N__47409\,
            I => \N__47399\
        );

    \I__11013\ : InMux
    port map (
            O => \N__47408\,
            I => \N__47396\
        );

    \I__11012\ : Odrv4
    port map (
            O => \N__47405\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__11011\ : Odrv12
    port map (
            O => \N__47402\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__11010\ : Odrv4
    port map (
            O => \N__47399\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__47396\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__11008\ : InMux
    port map (
            O => \N__47387\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__11007\ : CascadeMux
    port map (
            O => \N__47384\,
            I => \N__47380\
        );

    \I__11006\ : InMux
    port map (
            O => \N__47383\,
            I => \N__47377\
        );

    \I__11005\ : InMux
    port map (
            O => \N__47380\,
            I => \N__47374\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__47377\,
            I => \N__47371\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__47374\,
            I => \N__47368\
        );

    \I__11002\ : Span4Mux_h
    port map (
            O => \N__47371\,
            I => \N__47363\
        );

    \I__11001\ : Span4Mux_v
    port map (
            O => \N__47368\,
            I => \N__47360\
        );

    \I__11000\ : InMux
    port map (
            O => \N__47367\,
            I => \N__47355\
        );

    \I__10999\ : InMux
    port map (
            O => \N__47366\,
            I => \N__47355\
        );

    \I__10998\ : Odrv4
    port map (
            O => \N__47363\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10997\ : Odrv4
    port map (
            O => \N__47360\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__47355\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10995\ : InMux
    port map (
            O => \N__47348\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__10994\ : CascadeMux
    port map (
            O => \N__47345\,
            I => \N__47342\
        );

    \I__10993\ : InMux
    port map (
            O => \N__47342\,
            I => \N__47337\
        );

    \I__10992\ : InMux
    port map (
            O => \N__47341\,
            I => \N__47334\
        );

    \I__10991\ : InMux
    port map (
            O => \N__47340\,
            I => \N__47331\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__47337\,
            I => \N__47328\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__47334\,
            I => \N__47323\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__47331\,
            I => \N__47323\
        );

    \I__10987\ : Span4Mux_v
    port map (
            O => \N__47328\,
            I => \N__47319\
        );

    \I__10986\ : Span4Mux_v
    port map (
            O => \N__47323\,
            I => \N__47316\
        );

    \I__10985\ : InMux
    port map (
            O => \N__47322\,
            I => \N__47313\
        );

    \I__10984\ : Odrv4
    port map (
            O => \N__47319\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10983\ : Odrv4
    port map (
            O => \N__47316\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__47313\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10981\ : InMux
    port map (
            O => \N__47306\,
            I => \N__47302\
        );

    \I__10980\ : CascadeMux
    port map (
            O => \N__47305\,
            I => \N__47298\
        );

    \I__10979\ : LocalMux
    port map (
            O => \N__47302\,
            I => \N__47295\
        );

    \I__10978\ : InMux
    port map (
            O => \N__47301\,
            I => \N__47292\
        );

    \I__10977\ : InMux
    port map (
            O => \N__47298\,
            I => \N__47289\
        );

    \I__10976\ : Span4Mux_v
    port map (
            O => \N__47295\,
            I => \N__47284\
        );

    \I__10975\ : LocalMux
    port map (
            O => \N__47292\,
            I => \N__47284\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__47289\,
            I => \N__47278\
        );

    \I__10973\ : Span4Mux_v
    port map (
            O => \N__47284\,
            I => \N__47278\
        );

    \I__10972\ : InMux
    port map (
            O => \N__47283\,
            I => \N__47275\
        );

    \I__10971\ : Span4Mux_h
    port map (
            O => \N__47278\,
            I => \N__47272\
        );

    \I__10970\ : LocalMux
    port map (
            O => \N__47275\,
            I => \N__47269\
        );

    \I__10969\ : Odrv4
    port map (
            O => \N__47272\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__10968\ : Odrv4
    port map (
            O => \N__47269\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__10967\ : InMux
    port map (
            O => \N__47264\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__10966\ : CascadeMux
    port map (
            O => \N__47261\,
            I => \N__47257\
        );

    \I__10965\ : InMux
    port map (
            O => \N__47260\,
            I => \N__47252\
        );

    \I__10964\ : InMux
    port map (
            O => \N__47257\,
            I => \N__47249\
        );

    \I__10963\ : InMux
    port map (
            O => \N__47256\,
            I => \N__47244\
        );

    \I__10962\ : InMux
    port map (
            O => \N__47255\,
            I => \N__47244\
        );

    \I__10961\ : LocalMux
    port map (
            O => \N__47252\,
            I => \N__47241\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__47249\,
            I => \N__47238\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__47244\,
            I => \N__47235\
        );

    \I__10958\ : Span4Mux_h
    port map (
            O => \N__47241\,
            I => \N__47232\
        );

    \I__10957\ : Span4Mux_v
    port map (
            O => \N__47238\,
            I => \N__47227\
        );

    \I__10956\ : Span4Mux_h
    port map (
            O => \N__47235\,
            I => \N__47227\
        );

    \I__10955\ : Odrv4
    port map (
            O => \N__47232\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__10954\ : Odrv4
    port map (
            O => \N__47227\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__10953\ : InMux
    port map (
            O => \N__47222\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__10952\ : InMux
    port map (
            O => \N__47219\,
            I => \N__47212\
        );

    \I__10951\ : InMux
    port map (
            O => \N__47218\,
            I => \N__47212\
        );

    \I__10950\ : InMux
    port map (
            O => \N__47217\,
            I => \N__47209\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__47212\,
            I => \N__47204\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__47209\,
            I => \N__47204\
        );

    \I__10947\ : Span4Mux_h
    port map (
            O => \N__47204\,
            I => \N__47201\
        );

    \I__10946\ : Span4Mux_v
    port map (
            O => \N__47201\,
            I => \N__47197\
        );

    \I__10945\ : InMux
    port map (
            O => \N__47200\,
            I => \N__47194\
        );

    \I__10944\ : Odrv4
    port map (
            O => \N__47197\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__47194\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__10942\ : InMux
    port map (
            O => \N__47189\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__10941\ : CascadeMux
    port map (
            O => \N__47186\,
            I => \N__47183\
        );

    \I__10940\ : InMux
    port map (
            O => \N__47183\,
            I => \N__47180\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__47180\,
            I => \N__47175\
        );

    \I__10938\ : InMux
    port map (
            O => \N__47179\,
            I => \N__47172\
        );

    \I__10937\ : InMux
    port map (
            O => \N__47178\,
            I => \N__47169\
        );

    \I__10936\ : Span4Mux_h
    port map (
            O => \N__47175\,
            I => \N__47164\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__47172\,
            I => \N__47164\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__47169\,
            I => \N__47160\
        );

    \I__10933\ : Span4Mux_v
    port map (
            O => \N__47164\,
            I => \N__47157\
        );

    \I__10932\ : InMux
    port map (
            O => \N__47163\,
            I => \N__47154\
        );

    \I__10931\ : Odrv12
    port map (
            O => \N__47160\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10930\ : Odrv4
    port map (
            O => \N__47157\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10929\ : LocalMux
    port map (
            O => \N__47154\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10928\ : InMux
    port map (
            O => \N__47147\,
            I => \bfn_18_20_0_\
        );

    \I__10927\ : CascadeMux
    port map (
            O => \N__47144\,
            I => \N__47141\
        );

    \I__10926\ : InMux
    port map (
            O => \N__47141\,
            I => \N__47137\
        );

    \I__10925\ : InMux
    port map (
            O => \N__47140\,
            I => \N__47134\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__47137\,
            I => \N__47131\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__47134\,
            I => \N__47126\
        );

    \I__10922\ : Span4Mux_h
    port map (
            O => \N__47131\,
            I => \N__47123\
        );

    \I__10921\ : InMux
    port map (
            O => \N__47130\,
            I => \N__47118\
        );

    \I__10920\ : InMux
    port map (
            O => \N__47129\,
            I => \N__47118\
        );

    \I__10919\ : Span4Mux_h
    port map (
            O => \N__47126\,
            I => \N__47113\
        );

    \I__10918\ : Span4Mux_v
    port map (
            O => \N__47123\,
            I => \N__47113\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__47118\,
            I => \N__47110\
        );

    \I__10916\ : Odrv4
    port map (
            O => \N__47113\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10915\ : Odrv12
    port map (
            O => \N__47110\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10914\ : InMux
    port map (
            O => \N__47105\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__10913\ : CascadeMux
    port map (
            O => \N__47102\,
            I => \N__47099\
        );

    \I__10912\ : InMux
    port map (
            O => \N__47099\,
            I => \N__47095\
        );

    \I__10911\ : InMux
    port map (
            O => \N__47098\,
            I => \N__47092\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__47095\,
            I => \N__47085\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__47092\,
            I => \N__47085\
        );

    \I__10908\ : InMux
    port map (
            O => \N__47091\,
            I => \N__47082\
        );

    \I__10907\ : InMux
    port map (
            O => \N__47090\,
            I => \N__47079\
        );

    \I__10906\ : Span4Mux_v
    port map (
            O => \N__47085\,
            I => \N__47076\
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__47082\,
            I => \N__47073\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__47079\,
            I => \N__47070\
        );

    \I__10903\ : Odrv4
    port map (
            O => \N__47076\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10902\ : Odrv12
    port map (
            O => \N__47073\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10901\ : Odrv4
    port map (
            O => \N__47070\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10900\ : InMux
    port map (
            O => \N__47063\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__10899\ : CascadeMux
    port map (
            O => \N__47060\,
            I => \N__47057\
        );

    \I__10898\ : InMux
    port map (
            O => \N__47057\,
            I => \N__47053\
        );

    \I__10897\ : CascadeMux
    port map (
            O => \N__47056\,
            I => \N__47050\
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__47053\,
            I => \N__47045\
        );

    \I__10895\ : InMux
    port map (
            O => \N__47050\,
            I => \N__47042\
        );

    \I__10894\ : InMux
    port map (
            O => \N__47049\,
            I => \N__47039\
        );

    \I__10893\ : InMux
    port map (
            O => \N__47048\,
            I => \N__47036\
        );

    \I__10892\ : Span4Mux_h
    port map (
            O => \N__47045\,
            I => \N__47033\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__47042\,
            I => \N__47028\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__47039\,
            I => \N__47028\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__47036\,
            I => \N__47025\
        );

    \I__10888\ : Span4Mux_v
    port map (
            O => \N__47033\,
            I => \N__47020\
        );

    \I__10887\ : Span4Mux_h
    port map (
            O => \N__47028\,
            I => \N__47020\
        );

    \I__10886\ : Odrv12
    port map (
            O => \N__47025\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10885\ : Odrv4
    port map (
            O => \N__47020\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10884\ : InMux
    port map (
            O => \N__47015\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__10883\ : InMux
    port map (
            O => \N__47012\,
            I => \N__47008\
        );

    \I__10882\ : InMux
    port map (
            O => \N__47011\,
            I => \N__47004\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__47008\,
            I => \N__47000\
        );

    \I__10880\ : InMux
    port map (
            O => \N__47007\,
            I => \N__46997\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__47004\,
            I => \N__46994\
        );

    \I__10878\ : InMux
    port map (
            O => \N__47003\,
            I => \N__46991\
        );

    \I__10877\ : Span4Mux_v
    port map (
            O => \N__47000\,
            I => \N__46988\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__46997\,
            I => \N__46985\
        );

    \I__10875\ : Span4Mux_v
    port map (
            O => \N__46994\,
            I => \N__46980\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__46991\,
            I => \N__46980\
        );

    \I__10873\ : Odrv4
    port map (
            O => \N__46988\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10872\ : Odrv12
    port map (
            O => \N__46985\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10871\ : Odrv4
    port map (
            O => \N__46980\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10870\ : InMux
    port map (
            O => \N__46973\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__10869\ : InMux
    port map (
            O => \N__46970\,
            I => \N__46967\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__46967\,
            I => \N__46964\
        );

    \I__10867\ : Span4Mux_v
    port map (
            O => \N__46964\,
            I => \N__46961\
        );

    \I__10866\ : Odrv4
    port map (
            O => \N__46961\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__10865\ : InMux
    port map (
            O => \N__46958\,
            I => \N__46955\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__46955\,
            I => \N__46952\
        );

    \I__10863\ : Odrv4
    port map (
            O => \N__46952\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__10862\ : InMux
    port map (
            O => \N__46949\,
            I => \N__46946\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__46946\,
            I => \N__46943\
        );

    \I__10860\ : Odrv4
    port map (
            O => \N__46943\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__10859\ : InMux
    port map (
            O => \N__46940\,
            I => \N__46937\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__46937\,
            I => \N__46934\
        );

    \I__10857\ : Odrv4
    port map (
            O => \N__46934\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__10856\ : CascadeMux
    port map (
            O => \N__46931\,
            I => \N__46927\
        );

    \I__10855\ : CascadeMux
    port map (
            O => \N__46930\,
            I => \N__46924\
        );

    \I__10854\ : InMux
    port map (
            O => \N__46927\,
            I => \N__46921\
        );

    \I__10853\ : InMux
    port map (
            O => \N__46924\,
            I => \N__46918\
        );

    \I__10852\ : LocalMux
    port map (
            O => \N__46921\,
            I => \N__46914\
        );

    \I__10851\ : LocalMux
    port map (
            O => \N__46918\,
            I => \N__46911\
        );

    \I__10850\ : InMux
    port map (
            O => \N__46917\,
            I => \N__46908\
        );

    \I__10849\ : Span4Mux_v
    port map (
            O => \N__46914\,
            I => \N__46905\
        );

    \I__10848\ : Span4Mux_v
    port map (
            O => \N__46911\,
            I => \N__46899\
        );

    \I__10847\ : LocalMux
    port map (
            O => \N__46908\,
            I => \N__46899\
        );

    \I__10846\ : Span4Mux_v
    port map (
            O => \N__46905\,
            I => \N__46896\
        );

    \I__10845\ : InMux
    port map (
            O => \N__46904\,
            I => \N__46893\
        );

    \I__10844\ : Span4Mux_h
    port map (
            O => \N__46899\,
            I => \N__46890\
        );

    \I__10843\ : Span4Mux_h
    port map (
            O => \N__46896\,
            I => \N__46885\
        );

    \I__10842\ : LocalMux
    port map (
            O => \N__46893\,
            I => \N__46885\
        );

    \I__10841\ : Odrv4
    port map (
            O => \N__46890\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10840\ : Odrv4
    port map (
            O => \N__46885\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10839\ : CascadeMux
    port map (
            O => \N__46880\,
            I => \N__46876\
        );

    \I__10838\ : CascadeMux
    port map (
            O => \N__46879\,
            I => \N__46873\
        );

    \I__10837\ : InMux
    port map (
            O => \N__46876\,
            I => \N__46868\
        );

    \I__10836\ : InMux
    port map (
            O => \N__46873\,
            I => \N__46868\
        );

    \I__10835\ : LocalMux
    port map (
            O => \N__46868\,
            I => \N__46864\
        );

    \I__10834\ : InMux
    port map (
            O => \N__46867\,
            I => \N__46861\
        );

    \I__10833\ : Span4Mux_v
    port map (
            O => \N__46864\,
            I => \N__46856\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__46861\,
            I => \N__46856\
        );

    \I__10831\ : Span4Mux_h
    port map (
            O => \N__46856\,
            I => \N__46852\
        );

    \I__10830\ : InMux
    port map (
            O => \N__46855\,
            I => \N__46849\
        );

    \I__10829\ : Odrv4
    port map (
            O => \N__46852\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__10828\ : LocalMux
    port map (
            O => \N__46849\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__10827\ : InMux
    port map (
            O => \N__46844\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__10826\ : CascadeMux
    port map (
            O => \N__46841\,
            I => \N__46837\
        );

    \I__10825\ : CascadeMux
    port map (
            O => \N__46840\,
            I => \N__46834\
        );

    \I__10824\ : InMux
    port map (
            O => \N__46837\,
            I => \N__46831\
        );

    \I__10823\ : InMux
    port map (
            O => \N__46834\,
            I => \N__46828\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__46831\,
            I => \N__46822\
        );

    \I__10821\ : LocalMux
    port map (
            O => \N__46828\,
            I => \N__46822\
        );

    \I__10820\ : InMux
    port map (
            O => \N__46827\,
            I => \N__46819\
        );

    \I__10819\ : Span4Mux_v
    port map (
            O => \N__46822\,
            I => \N__46815\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__46819\,
            I => \N__46812\
        );

    \I__10817\ : InMux
    port map (
            O => \N__46818\,
            I => \N__46809\
        );

    \I__10816\ : Span4Mux_v
    port map (
            O => \N__46815\,
            I => \N__46806\
        );

    \I__10815\ : Span4Mux_h
    port map (
            O => \N__46812\,
            I => \N__46801\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__46809\,
            I => \N__46801\
        );

    \I__10813\ : Odrv4
    port map (
            O => \N__46806\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__10812\ : Odrv4
    port map (
            O => \N__46801\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__10811\ : InMux
    port map (
            O => \N__46796\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__10810\ : CascadeMux
    port map (
            O => \N__46793\,
            I => \N__46790\
        );

    \I__10809\ : InMux
    port map (
            O => \N__46790\,
            I => \N__46786\
        );

    \I__10808\ : CascadeMux
    port map (
            O => \N__46789\,
            I => \N__46783\
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__46786\,
            I => \N__46778\
        );

    \I__10806\ : InMux
    port map (
            O => \N__46783\,
            I => \N__46775\
        );

    \I__10805\ : InMux
    port map (
            O => \N__46782\,
            I => \N__46772\
        );

    \I__10804\ : InMux
    port map (
            O => \N__46781\,
            I => \N__46769\
        );

    \I__10803\ : Span4Mux_v
    port map (
            O => \N__46778\,
            I => \N__46766\
        );

    \I__10802\ : LocalMux
    port map (
            O => \N__46775\,
            I => \N__46763\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__46772\,
            I => \N__46760\
        );

    \I__10800\ : LocalMux
    port map (
            O => \N__46769\,
            I => \N__46757\
        );

    \I__10799\ : Span4Mux_v
    port map (
            O => \N__46766\,
            I => \N__46754\
        );

    \I__10798\ : Span4Mux_v
    port map (
            O => \N__46763\,
            I => \N__46749\
        );

    \I__10797\ : Span4Mux_h
    port map (
            O => \N__46760\,
            I => \N__46749\
        );

    \I__10796\ : Span4Mux_v
    port map (
            O => \N__46757\,
            I => \N__46746\
        );

    \I__10795\ : Odrv4
    port map (
            O => \N__46754\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__10794\ : Odrv4
    port map (
            O => \N__46749\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__10793\ : Odrv4
    port map (
            O => \N__46746\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__10792\ : InMux
    port map (
            O => \N__46739\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__10791\ : InMux
    port map (
            O => \N__46736\,
            I => \N__46732\
        );

    \I__10790\ : InMux
    port map (
            O => \N__46735\,
            I => \N__46728\
        );

    \I__10789\ : LocalMux
    port map (
            O => \N__46732\,
            I => \N__46725\
        );

    \I__10788\ : InMux
    port map (
            O => \N__46731\,
            I => \N__46722\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__46728\,
            I => \N__46715\
        );

    \I__10786\ : Span4Mux_v
    port map (
            O => \N__46725\,
            I => \N__46715\
        );

    \I__10785\ : LocalMux
    port map (
            O => \N__46722\,
            I => \N__46715\
        );

    \I__10784\ : Span4Mux_v
    port map (
            O => \N__46715\,
            I => \N__46711\
        );

    \I__10783\ : InMux
    port map (
            O => \N__46714\,
            I => \N__46708\
        );

    \I__10782\ : Odrv4
    port map (
            O => \N__46711\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__46708\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10780\ : InMux
    port map (
            O => \N__46703\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__10779\ : CascadeMux
    port map (
            O => \N__46700\,
            I => \N__46696\
        );

    \I__10778\ : InMux
    port map (
            O => \N__46699\,
            I => \N__46693\
        );

    \I__10777\ : InMux
    port map (
            O => \N__46696\,
            I => \N__46690\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__46693\,
            I => \N__46687\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__46690\,
            I => \N__46681\
        );

    \I__10774\ : Span4Mux_h
    port map (
            O => \N__46687\,
            I => \N__46681\
        );

    \I__10773\ : InMux
    port map (
            O => \N__46686\,
            I => \N__46678\
        );

    \I__10772\ : Odrv4
    port map (
            O => \N__46681\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__46678\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__10770\ : CascadeMux
    port map (
            O => \N__46673\,
            I => \N__46670\
        );

    \I__10769\ : InMux
    port map (
            O => \N__46670\,
            I => \N__46667\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__46667\,
            I => \N__46664\
        );

    \I__10767\ : Odrv12
    port map (
            O => \N__46664\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\
        );

    \I__10766\ : CascadeMux
    port map (
            O => \N__46661\,
            I => \N__46654\
        );

    \I__10765\ : CascadeMux
    port map (
            O => \N__46660\,
            I => \N__46639\
        );

    \I__10764\ : CascadeMux
    port map (
            O => \N__46659\,
            I => \N__46633\
        );

    \I__10763\ : InMux
    port map (
            O => \N__46658\,
            I => \N__46614\
        );

    \I__10762\ : InMux
    port map (
            O => \N__46657\,
            I => \N__46614\
        );

    \I__10761\ : InMux
    port map (
            O => \N__46654\,
            I => \N__46614\
        );

    \I__10760\ : CascadeMux
    port map (
            O => \N__46653\,
            I => \N__46611\
        );

    \I__10759\ : CascadeMux
    port map (
            O => \N__46652\,
            I => \N__46607\
        );

    \I__10758\ : CascadeMux
    port map (
            O => \N__46651\,
            I => \N__46584\
        );

    \I__10757\ : InMux
    port map (
            O => \N__46650\,
            I => \N__46567\
        );

    \I__10756\ : InMux
    port map (
            O => \N__46649\,
            I => \N__46567\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46648\,
            I => \N__46567\
        );

    \I__10754\ : InMux
    port map (
            O => \N__46647\,
            I => \N__46567\
        );

    \I__10753\ : InMux
    port map (
            O => \N__46646\,
            I => \N__46567\
        );

    \I__10752\ : InMux
    port map (
            O => \N__46645\,
            I => \N__46567\
        );

    \I__10751\ : InMux
    port map (
            O => \N__46644\,
            I => \N__46567\
        );

    \I__10750\ : InMux
    port map (
            O => \N__46643\,
            I => \N__46567\
        );

    \I__10749\ : InMux
    port map (
            O => \N__46642\,
            I => \N__46543\
        );

    \I__10748\ : InMux
    port map (
            O => \N__46639\,
            I => \N__46543\
        );

    \I__10747\ : InMux
    port map (
            O => \N__46638\,
            I => \N__46543\
        );

    \I__10746\ : InMux
    port map (
            O => \N__46637\,
            I => \N__46543\
        );

    \I__10745\ : InMux
    port map (
            O => \N__46636\,
            I => \N__46543\
        );

    \I__10744\ : InMux
    port map (
            O => \N__46633\,
            I => \N__46543\
        );

    \I__10743\ : InMux
    port map (
            O => \N__46632\,
            I => \N__46543\
        );

    \I__10742\ : InMux
    port map (
            O => \N__46631\,
            I => \N__46543\
        );

    \I__10741\ : InMux
    port map (
            O => \N__46630\,
            I => \N__46528\
        );

    \I__10740\ : InMux
    port map (
            O => \N__46629\,
            I => \N__46528\
        );

    \I__10739\ : InMux
    port map (
            O => \N__46628\,
            I => \N__46528\
        );

    \I__10738\ : InMux
    port map (
            O => \N__46627\,
            I => \N__46528\
        );

    \I__10737\ : InMux
    port map (
            O => \N__46626\,
            I => \N__46528\
        );

    \I__10736\ : InMux
    port map (
            O => \N__46625\,
            I => \N__46528\
        );

    \I__10735\ : InMux
    port map (
            O => \N__46624\,
            I => \N__46528\
        );

    \I__10734\ : CascadeMux
    port map (
            O => \N__46623\,
            I => \N__46520\
        );

    \I__10733\ : CascadeMux
    port map (
            O => \N__46622\,
            I => \N__46517\
        );

    \I__10732\ : CascadeMux
    port map (
            O => \N__46621\,
            I => \N__46514\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__46614\,
            I => \N__46501\
        );

    \I__10730\ : InMux
    port map (
            O => \N__46611\,
            I => \N__46484\
        );

    \I__10729\ : InMux
    port map (
            O => \N__46610\,
            I => \N__46484\
        );

    \I__10728\ : InMux
    port map (
            O => \N__46607\,
            I => \N__46484\
        );

    \I__10727\ : InMux
    port map (
            O => \N__46606\,
            I => \N__46484\
        );

    \I__10726\ : InMux
    port map (
            O => \N__46605\,
            I => \N__46484\
        );

    \I__10725\ : InMux
    port map (
            O => \N__46604\,
            I => \N__46484\
        );

    \I__10724\ : InMux
    port map (
            O => \N__46603\,
            I => \N__46484\
        );

    \I__10723\ : InMux
    port map (
            O => \N__46602\,
            I => \N__46484\
        );

    \I__10722\ : InMux
    port map (
            O => \N__46601\,
            I => \N__46481\
        );

    \I__10721\ : CascadeMux
    port map (
            O => \N__46600\,
            I => \N__46478\
        );

    \I__10720\ : CascadeMux
    port map (
            O => \N__46599\,
            I => \N__46474\
        );

    \I__10719\ : CascadeMux
    port map (
            O => \N__46598\,
            I => \N__46470\
        );

    \I__10718\ : CascadeMux
    port map (
            O => \N__46597\,
            I => \N__46466\
        );

    \I__10717\ : CascadeMux
    port map (
            O => \N__46596\,
            I => \N__46463\
        );

    \I__10716\ : CascadeMux
    port map (
            O => \N__46595\,
            I => \N__46459\
        );

    \I__10715\ : CascadeMux
    port map (
            O => \N__46594\,
            I => \N__46455\
        );

    \I__10714\ : CascadeMux
    port map (
            O => \N__46593\,
            I => \N__46451\
        );

    \I__10713\ : CascadeMux
    port map (
            O => \N__46592\,
            I => \N__46435\
        );

    \I__10712\ : CascadeMux
    port map (
            O => \N__46591\,
            I => \N__46431\
        );

    \I__10711\ : CascadeMux
    port map (
            O => \N__46590\,
            I => \N__46427\
        );

    \I__10710\ : InMux
    port map (
            O => \N__46589\,
            I => \N__46420\
        );

    \I__10709\ : InMux
    port map (
            O => \N__46588\,
            I => \N__46420\
        );

    \I__10708\ : InMux
    port map (
            O => \N__46587\,
            I => \N__46420\
        );

    \I__10707\ : InMux
    port map (
            O => \N__46584\,
            I => \N__46417\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__46567\,
            I => \N__46414\
        );

    \I__10705\ : InMux
    port map (
            O => \N__46566\,
            I => \N__46399\
        );

    \I__10704\ : InMux
    port map (
            O => \N__46565\,
            I => \N__46399\
        );

    \I__10703\ : InMux
    port map (
            O => \N__46564\,
            I => \N__46399\
        );

    \I__10702\ : InMux
    port map (
            O => \N__46563\,
            I => \N__46399\
        );

    \I__10701\ : InMux
    port map (
            O => \N__46562\,
            I => \N__46399\
        );

    \I__10700\ : InMux
    port map (
            O => \N__46561\,
            I => \N__46399\
        );

    \I__10699\ : InMux
    port map (
            O => \N__46560\,
            I => \N__46399\
        );

    \I__10698\ : LocalMux
    port map (
            O => \N__46543\,
            I => \N__46394\
        );

    \I__10697\ : LocalMux
    port map (
            O => \N__46528\,
            I => \N__46394\
        );

    \I__10696\ : InMux
    port map (
            O => \N__46527\,
            I => \N__46389\
        );

    \I__10695\ : InMux
    port map (
            O => \N__46526\,
            I => \N__46389\
        );

    \I__10694\ : InMux
    port map (
            O => \N__46525\,
            I => \N__46378\
        );

    \I__10693\ : InMux
    port map (
            O => \N__46524\,
            I => \N__46378\
        );

    \I__10692\ : InMux
    port map (
            O => \N__46523\,
            I => \N__46378\
        );

    \I__10691\ : InMux
    port map (
            O => \N__46520\,
            I => \N__46378\
        );

    \I__10690\ : InMux
    port map (
            O => \N__46517\,
            I => \N__46378\
        );

    \I__10689\ : InMux
    port map (
            O => \N__46514\,
            I => \N__46368\
        );

    \I__10688\ : InMux
    port map (
            O => \N__46513\,
            I => \N__46368\
        );

    \I__10687\ : InMux
    port map (
            O => \N__46512\,
            I => \N__46368\
        );

    \I__10686\ : CascadeMux
    port map (
            O => \N__46511\,
            I => \N__46364\
        );

    \I__10685\ : CascadeMux
    port map (
            O => \N__46510\,
            I => \N__46360\
        );

    \I__10684\ : CascadeMux
    port map (
            O => \N__46509\,
            I => \N__46356\
        );

    \I__10683\ : CascadeMux
    port map (
            O => \N__46508\,
            I => \N__46352\
        );

    \I__10682\ : CascadeMux
    port map (
            O => \N__46507\,
            I => \N__46349\
        );

    \I__10681\ : CascadeMux
    port map (
            O => \N__46506\,
            I => \N__46345\
        );

    \I__10680\ : CascadeMux
    port map (
            O => \N__46505\,
            I => \N__46341\
        );

    \I__10679\ : CascadeMux
    port map (
            O => \N__46504\,
            I => \N__46337\
        );

    \I__10678\ : Span4Mux_v
    port map (
            O => \N__46501\,
            I => \N__46333\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__46484\,
            I => \N__46328\
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__46481\,
            I => \N__46328\
        );

    \I__10675\ : InMux
    port map (
            O => \N__46478\,
            I => \N__46313\
        );

    \I__10674\ : InMux
    port map (
            O => \N__46477\,
            I => \N__46313\
        );

    \I__10673\ : InMux
    port map (
            O => \N__46474\,
            I => \N__46313\
        );

    \I__10672\ : InMux
    port map (
            O => \N__46473\,
            I => \N__46313\
        );

    \I__10671\ : InMux
    port map (
            O => \N__46470\,
            I => \N__46313\
        );

    \I__10670\ : InMux
    port map (
            O => \N__46469\,
            I => \N__46313\
        );

    \I__10669\ : InMux
    port map (
            O => \N__46466\,
            I => \N__46313\
        );

    \I__10668\ : InMux
    port map (
            O => \N__46463\,
            I => \N__46296\
        );

    \I__10667\ : InMux
    port map (
            O => \N__46462\,
            I => \N__46296\
        );

    \I__10666\ : InMux
    port map (
            O => \N__46459\,
            I => \N__46296\
        );

    \I__10665\ : InMux
    port map (
            O => \N__46458\,
            I => \N__46296\
        );

    \I__10664\ : InMux
    port map (
            O => \N__46455\,
            I => \N__46296\
        );

    \I__10663\ : InMux
    port map (
            O => \N__46454\,
            I => \N__46296\
        );

    \I__10662\ : InMux
    port map (
            O => \N__46451\,
            I => \N__46296\
        );

    \I__10661\ : InMux
    port map (
            O => \N__46450\,
            I => \N__46296\
        );

    \I__10660\ : CascadeMux
    port map (
            O => \N__46449\,
            I => \N__46293\
        );

    \I__10659\ : CascadeMux
    port map (
            O => \N__46448\,
            I => \N__46289\
        );

    \I__10658\ : CascadeMux
    port map (
            O => \N__46447\,
            I => \N__46285\
        );

    \I__10657\ : CascadeMux
    port map (
            O => \N__46446\,
            I => \N__46281\
        );

    \I__10656\ : CascadeMux
    port map (
            O => \N__46445\,
            I => \N__46277\
        );

    \I__10655\ : CascadeMux
    port map (
            O => \N__46444\,
            I => \N__46273\
        );

    \I__10654\ : CascadeMux
    port map (
            O => \N__46443\,
            I => \N__46269\
        );

    \I__10653\ : CascadeMux
    port map (
            O => \N__46442\,
            I => \N__46265\
        );

    \I__10652\ : CascadeMux
    port map (
            O => \N__46441\,
            I => \N__46261\
        );

    \I__10651\ : CascadeMux
    port map (
            O => \N__46440\,
            I => \N__46257\
        );

    \I__10650\ : CascadeMux
    port map (
            O => \N__46439\,
            I => \N__46253\
        );

    \I__10649\ : InMux
    port map (
            O => \N__46438\,
            I => \N__46239\
        );

    \I__10648\ : InMux
    port map (
            O => \N__46435\,
            I => \N__46239\
        );

    \I__10647\ : InMux
    port map (
            O => \N__46434\,
            I => \N__46239\
        );

    \I__10646\ : InMux
    port map (
            O => \N__46431\,
            I => \N__46239\
        );

    \I__10645\ : InMux
    port map (
            O => \N__46430\,
            I => \N__46239\
        );

    \I__10644\ : InMux
    port map (
            O => \N__46427\,
            I => \N__46239\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__46420\,
            I => \N__46236\
        );

    \I__10642\ : LocalMux
    port map (
            O => \N__46417\,
            I => \N__46229\
        );

    \I__10641\ : Span12Mux_s11_h
    port map (
            O => \N__46414\,
            I => \N__46229\
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__46399\,
            I => \N__46229\
        );

    \I__10639\ : Span4Mux_v
    port map (
            O => \N__46394\,
            I => \N__46222\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__46389\,
            I => \N__46222\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__46378\,
            I => \N__46222\
        );

    \I__10636\ : InMux
    port map (
            O => \N__46377\,
            I => \N__46215\
        );

    \I__10635\ : InMux
    port map (
            O => \N__46376\,
            I => \N__46215\
        );

    \I__10634\ : InMux
    port map (
            O => \N__46375\,
            I => \N__46215\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__46368\,
            I => \N__46212\
        );

    \I__10632\ : InMux
    port map (
            O => \N__46367\,
            I => \N__46195\
        );

    \I__10631\ : InMux
    port map (
            O => \N__46364\,
            I => \N__46195\
        );

    \I__10630\ : InMux
    port map (
            O => \N__46363\,
            I => \N__46195\
        );

    \I__10629\ : InMux
    port map (
            O => \N__46360\,
            I => \N__46195\
        );

    \I__10628\ : InMux
    port map (
            O => \N__46359\,
            I => \N__46195\
        );

    \I__10627\ : InMux
    port map (
            O => \N__46356\,
            I => \N__46195\
        );

    \I__10626\ : InMux
    port map (
            O => \N__46355\,
            I => \N__46195\
        );

    \I__10625\ : InMux
    port map (
            O => \N__46352\,
            I => \N__46195\
        );

    \I__10624\ : InMux
    port map (
            O => \N__46349\,
            I => \N__46178\
        );

    \I__10623\ : InMux
    port map (
            O => \N__46348\,
            I => \N__46178\
        );

    \I__10622\ : InMux
    port map (
            O => \N__46345\,
            I => \N__46178\
        );

    \I__10621\ : InMux
    port map (
            O => \N__46344\,
            I => \N__46178\
        );

    \I__10620\ : InMux
    port map (
            O => \N__46341\,
            I => \N__46178\
        );

    \I__10619\ : InMux
    port map (
            O => \N__46340\,
            I => \N__46178\
        );

    \I__10618\ : InMux
    port map (
            O => \N__46337\,
            I => \N__46178\
        );

    \I__10617\ : InMux
    port map (
            O => \N__46336\,
            I => \N__46178\
        );

    \I__10616\ : Span4Mux_h
    port map (
            O => \N__46333\,
            I => \N__46169\
        );

    \I__10615\ : Span4Mux_h
    port map (
            O => \N__46328\,
            I => \N__46169\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__46313\,
            I => \N__46169\
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__46296\,
            I => \N__46169\
        );

    \I__10612\ : InMux
    port map (
            O => \N__46293\,
            I => \N__46152\
        );

    \I__10611\ : InMux
    port map (
            O => \N__46292\,
            I => \N__46152\
        );

    \I__10610\ : InMux
    port map (
            O => \N__46289\,
            I => \N__46152\
        );

    \I__10609\ : InMux
    port map (
            O => \N__46288\,
            I => \N__46152\
        );

    \I__10608\ : InMux
    port map (
            O => \N__46285\,
            I => \N__46152\
        );

    \I__10607\ : InMux
    port map (
            O => \N__46284\,
            I => \N__46152\
        );

    \I__10606\ : InMux
    port map (
            O => \N__46281\,
            I => \N__46152\
        );

    \I__10605\ : InMux
    port map (
            O => \N__46280\,
            I => \N__46152\
        );

    \I__10604\ : InMux
    port map (
            O => \N__46277\,
            I => \N__46135\
        );

    \I__10603\ : InMux
    port map (
            O => \N__46276\,
            I => \N__46135\
        );

    \I__10602\ : InMux
    port map (
            O => \N__46273\,
            I => \N__46135\
        );

    \I__10601\ : InMux
    port map (
            O => \N__46272\,
            I => \N__46135\
        );

    \I__10600\ : InMux
    port map (
            O => \N__46269\,
            I => \N__46135\
        );

    \I__10599\ : InMux
    port map (
            O => \N__46268\,
            I => \N__46135\
        );

    \I__10598\ : InMux
    port map (
            O => \N__46265\,
            I => \N__46135\
        );

    \I__10597\ : InMux
    port map (
            O => \N__46264\,
            I => \N__46135\
        );

    \I__10596\ : InMux
    port map (
            O => \N__46261\,
            I => \N__46122\
        );

    \I__10595\ : InMux
    port map (
            O => \N__46260\,
            I => \N__46122\
        );

    \I__10594\ : InMux
    port map (
            O => \N__46257\,
            I => \N__46122\
        );

    \I__10593\ : InMux
    port map (
            O => \N__46256\,
            I => \N__46122\
        );

    \I__10592\ : InMux
    port map (
            O => \N__46253\,
            I => \N__46122\
        );

    \I__10591\ : InMux
    port map (
            O => \N__46252\,
            I => \N__46122\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__46239\,
            I => \N__46119\
        );

    \I__10589\ : Odrv12
    port map (
            O => \N__46236\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10588\ : Odrv12
    port map (
            O => \N__46229\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10587\ : Odrv4
    port map (
            O => \N__46222\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__46215\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10585\ : Odrv4
    port map (
            O => \N__46212\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__46195\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__46178\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10582\ : Odrv4
    port map (
            O => \N__46169\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__46152\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__46135\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__46122\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10578\ : Odrv4
    port map (
            O => \N__46119\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10577\ : InMux
    port map (
            O => \N__46094\,
            I => \N__46089\
        );

    \I__10576\ : InMux
    port map (
            O => \N__46093\,
            I => \N__46086\
        );

    \I__10575\ : InMux
    port map (
            O => \N__46092\,
            I => \N__46083\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__46089\,
            I => \N__46080\
        );

    \I__10573\ : LocalMux
    port map (
            O => \N__46086\,
            I => \N__46077\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__46083\,
            I => \N__46074\
        );

    \I__10571\ : Span4Mux_h
    port map (
            O => \N__46080\,
            I => \N__46071\
        );

    \I__10570\ : Span4Mux_h
    port map (
            O => \N__46077\,
            I => \N__46068\
        );

    \I__10569\ : Span4Mux_h
    port map (
            O => \N__46074\,
            I => \N__46065\
        );

    \I__10568\ : Odrv4
    port map (
            O => \N__46071\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10567\ : Odrv4
    port map (
            O => \N__46068\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10566\ : Odrv4
    port map (
            O => \N__46065\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10565\ : CascadeMux
    port map (
            O => \N__46058\,
            I => \N__46055\
        );

    \I__10564\ : InMux
    port map (
            O => \N__46055\,
            I => \N__46052\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__46052\,
            I => \N__46049\
        );

    \I__10562\ : Odrv12
    port map (
            O => \N__46049\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\
        );

    \I__10561\ : InMux
    port map (
            O => \N__46046\,
            I => \N__46042\
        );

    \I__10560\ : InMux
    port map (
            O => \N__46045\,
            I => \N__46038\
        );

    \I__10559\ : LocalMux
    port map (
            O => \N__46042\,
            I => \N__46035\
        );

    \I__10558\ : InMux
    port map (
            O => \N__46041\,
            I => \N__46032\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__46038\,
            I => \N__46029\
        );

    \I__10556\ : Span4Mux_h
    port map (
            O => \N__46035\,
            I => \N__46026\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__46032\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10554\ : Odrv12
    port map (
            O => \N__46029\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10553\ : Odrv4
    port map (
            O => \N__46026\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10552\ : CascadeMux
    port map (
            O => \N__46019\,
            I => \N__46016\
        );

    \I__10551\ : InMux
    port map (
            O => \N__46016\,
            I => \N__46013\
        );

    \I__10550\ : LocalMux
    port map (
            O => \N__46013\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__10549\ : InMux
    port map (
            O => \N__46010\,
            I => \N__45996\
        );

    \I__10548\ : CascadeMux
    port map (
            O => \N__46009\,
            I => \N__45988\
        );

    \I__10547\ : InMux
    port map (
            O => \N__46008\,
            I => \N__45975\
        );

    \I__10546\ : InMux
    port map (
            O => \N__46007\,
            I => \N__45975\
        );

    \I__10545\ : InMux
    port map (
            O => \N__46006\,
            I => \N__45975\
        );

    \I__10544\ : InMux
    port map (
            O => \N__46005\,
            I => \N__45975\
        );

    \I__10543\ : InMux
    port map (
            O => \N__46004\,
            I => \N__45966\
        );

    \I__10542\ : InMux
    port map (
            O => \N__46003\,
            I => \N__45966\
        );

    \I__10541\ : InMux
    port map (
            O => \N__46002\,
            I => \N__45966\
        );

    \I__10540\ : InMux
    port map (
            O => \N__46001\,
            I => \N__45966\
        );

    \I__10539\ : InMux
    port map (
            O => \N__46000\,
            I => \N__45963\
        );

    \I__10538\ : InMux
    port map (
            O => \N__45999\,
            I => \N__45952\
        );

    \I__10537\ : LocalMux
    port map (
            O => \N__45996\,
            I => \N__45949\
        );

    \I__10536\ : InMux
    port map (
            O => \N__45995\,
            I => \N__45944\
        );

    \I__10535\ : InMux
    port map (
            O => \N__45994\,
            I => \N__45944\
        );

    \I__10534\ : InMux
    port map (
            O => \N__45993\,
            I => \N__45937\
        );

    \I__10533\ : InMux
    port map (
            O => \N__45992\,
            I => \N__45937\
        );

    \I__10532\ : InMux
    port map (
            O => \N__45991\,
            I => \N__45937\
        );

    \I__10531\ : InMux
    port map (
            O => \N__45988\,
            I => \N__45926\
        );

    \I__10530\ : InMux
    port map (
            O => \N__45987\,
            I => \N__45926\
        );

    \I__10529\ : InMux
    port map (
            O => \N__45986\,
            I => \N__45926\
        );

    \I__10528\ : InMux
    port map (
            O => \N__45985\,
            I => \N__45926\
        );

    \I__10527\ : InMux
    port map (
            O => \N__45984\,
            I => \N__45926\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__45975\,
            I => \N__45919\
        );

    \I__10525\ : LocalMux
    port map (
            O => \N__45966\,
            I => \N__45919\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__45963\,
            I => \N__45919\
        );

    \I__10523\ : InMux
    port map (
            O => \N__45962\,
            I => \N__45900\
        );

    \I__10522\ : InMux
    port map (
            O => \N__45961\,
            I => \N__45900\
        );

    \I__10521\ : InMux
    port map (
            O => \N__45960\,
            I => \N__45900\
        );

    \I__10520\ : InMux
    port map (
            O => \N__45959\,
            I => \N__45891\
        );

    \I__10519\ : InMux
    port map (
            O => \N__45958\,
            I => \N__45891\
        );

    \I__10518\ : InMux
    port map (
            O => \N__45957\,
            I => \N__45891\
        );

    \I__10517\ : InMux
    port map (
            O => \N__45956\,
            I => \N__45891\
        );

    \I__10516\ : InMux
    port map (
            O => \N__45955\,
            I => \N__45888\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__45952\,
            I => \N__45856\
        );

    \I__10514\ : Span4Mux_h
    port map (
            O => \N__45949\,
            I => \N__45856\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__45944\,
            I => \N__45856\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__45937\,
            I => \N__45856\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__45926\,
            I => \N__45856\
        );

    \I__10510\ : Span4Mux_v
    port map (
            O => \N__45919\,
            I => \N__45856\
        );

    \I__10509\ : InMux
    port map (
            O => \N__45918\,
            I => \N__45839\
        );

    \I__10508\ : InMux
    port map (
            O => \N__45917\,
            I => \N__45839\
        );

    \I__10507\ : InMux
    port map (
            O => \N__45916\,
            I => \N__45839\
        );

    \I__10506\ : InMux
    port map (
            O => \N__45915\,
            I => \N__45839\
        );

    \I__10505\ : InMux
    port map (
            O => \N__45914\,
            I => \N__45839\
        );

    \I__10504\ : InMux
    port map (
            O => \N__45913\,
            I => \N__45839\
        );

    \I__10503\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45839\
        );

    \I__10502\ : InMux
    port map (
            O => \N__45911\,
            I => \N__45839\
        );

    \I__10501\ : CascadeMux
    port map (
            O => \N__45910\,
            I => \N__45827\
        );

    \I__10500\ : InMux
    port map (
            O => \N__45909\,
            I => \N__45819\
        );

    \I__10499\ : InMux
    port map (
            O => \N__45908\,
            I => \N__45819\
        );

    \I__10498\ : InMux
    port map (
            O => \N__45907\,
            I => \N__45819\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__45900\,
            I => \N__45814\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__45891\,
            I => \N__45814\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__45888\,
            I => \N__45810\
        );

    \I__10494\ : InMux
    port map (
            O => \N__45887\,
            I => \N__45795\
        );

    \I__10493\ : InMux
    port map (
            O => \N__45886\,
            I => \N__45795\
        );

    \I__10492\ : InMux
    port map (
            O => \N__45885\,
            I => \N__45795\
        );

    \I__10491\ : InMux
    port map (
            O => \N__45884\,
            I => \N__45795\
        );

    \I__10490\ : InMux
    port map (
            O => \N__45883\,
            I => \N__45795\
        );

    \I__10489\ : InMux
    port map (
            O => \N__45882\,
            I => \N__45795\
        );

    \I__10488\ : InMux
    port map (
            O => \N__45881\,
            I => \N__45795\
        );

    \I__10487\ : InMux
    port map (
            O => \N__45880\,
            I => \N__45780\
        );

    \I__10486\ : InMux
    port map (
            O => \N__45879\,
            I => \N__45780\
        );

    \I__10485\ : InMux
    port map (
            O => \N__45878\,
            I => \N__45780\
        );

    \I__10484\ : InMux
    port map (
            O => \N__45877\,
            I => \N__45780\
        );

    \I__10483\ : InMux
    port map (
            O => \N__45876\,
            I => \N__45780\
        );

    \I__10482\ : InMux
    port map (
            O => \N__45875\,
            I => \N__45780\
        );

    \I__10481\ : InMux
    port map (
            O => \N__45874\,
            I => \N__45780\
        );

    \I__10480\ : InMux
    port map (
            O => \N__45873\,
            I => \N__45775\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45872\,
            I => \N__45775\
        );

    \I__10478\ : InMux
    port map (
            O => \N__45871\,
            I => \N__45768\
        );

    \I__10477\ : InMux
    port map (
            O => \N__45870\,
            I => \N__45768\
        );

    \I__10476\ : InMux
    port map (
            O => \N__45869\,
            I => \N__45768\
        );

    \I__10475\ : Span4Mux_v
    port map (
            O => \N__45856\,
            I => \N__45763\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__45839\,
            I => \N__45763\
        );

    \I__10473\ : InMux
    port map (
            O => \N__45838\,
            I => \N__45752\
        );

    \I__10472\ : InMux
    port map (
            O => \N__45837\,
            I => \N__45752\
        );

    \I__10471\ : InMux
    port map (
            O => \N__45836\,
            I => \N__45752\
        );

    \I__10470\ : InMux
    port map (
            O => \N__45835\,
            I => \N__45752\
        );

    \I__10469\ : InMux
    port map (
            O => \N__45834\,
            I => \N__45752\
        );

    \I__10468\ : InMux
    port map (
            O => \N__45833\,
            I => \N__45745\
        );

    \I__10467\ : InMux
    port map (
            O => \N__45832\,
            I => \N__45745\
        );

    \I__10466\ : InMux
    port map (
            O => \N__45831\,
            I => \N__45745\
        );

    \I__10465\ : InMux
    port map (
            O => \N__45830\,
            I => \N__45738\
        );

    \I__10464\ : InMux
    port map (
            O => \N__45827\,
            I => \N__45738\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45826\,
            I => \N__45738\
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__45819\,
            I => \N__45733\
        );

    \I__10461\ : Span4Mux_v
    port map (
            O => \N__45814\,
            I => \N__45733\
        );

    \I__10460\ : InMux
    port map (
            O => \N__45813\,
            I => \N__45730\
        );

    \I__10459\ : Span12Mux_s11_v
    port map (
            O => \N__45810\,
            I => \N__45719\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__45795\,
            I => \N__45719\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__45780\,
            I => \N__45719\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__45775\,
            I => \N__45719\
        );

    \I__10455\ : LocalMux
    port map (
            O => \N__45768\,
            I => \N__45719\
        );

    \I__10454\ : Span4Mux_v
    port map (
            O => \N__45763\,
            I => \N__45716\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__45752\,
            I => \N__45705\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__45745\,
            I => \N__45705\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__45738\,
            I => \N__45705\
        );

    \I__10450\ : Sp12to4
    port map (
            O => \N__45733\,
            I => \N__45705\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__45730\,
            I => \N__45705\
        );

    \I__10448\ : Span12Mux_s11_h
    port map (
            O => \N__45719\,
            I => \N__45702\
        );

    \I__10447\ : Odrv4
    port map (
            O => \N__45716\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10446\ : Odrv12
    port map (
            O => \N__45705\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10445\ : Odrv12
    port map (
            O => \N__45702\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10444\ : InMux
    port map (
            O => \N__45695\,
            I => \N__45692\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__45692\,
            I => \N__45689\
        );

    \I__10442\ : Odrv4
    port map (
            O => \N__45689\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__10441\ : InMux
    port map (
            O => \N__45686\,
            I => \N__45682\
        );

    \I__10440\ : InMux
    port map (
            O => \N__45685\,
            I => \N__45679\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__45682\,
            I => \N__45676\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__45679\,
            I => \N__45673\
        );

    \I__10437\ : Span4Mux_h
    port map (
            O => \N__45676\,
            I => \N__45668\
        );

    \I__10436\ : Span4Mux_h
    port map (
            O => \N__45673\,
            I => \N__45665\
        );

    \I__10435\ : InMux
    port map (
            O => \N__45672\,
            I => \N__45660\
        );

    \I__10434\ : InMux
    port map (
            O => \N__45671\,
            I => \N__45660\
        );

    \I__10433\ : Odrv4
    port map (
            O => \N__45668\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__10432\ : Odrv4
    port map (
            O => \N__45665\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__45660\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__10430\ : CascadeMux
    port map (
            O => \N__45653\,
            I => \N__45650\
        );

    \I__10429\ : InMux
    port map (
            O => \N__45650\,
            I => \N__45647\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__45647\,
            I => \N__45644\
        );

    \I__10427\ : Span4Mux_h
    port map (
            O => \N__45644\,
            I => \N__45641\
        );

    \I__10426\ : Odrv4
    port map (
            O => \N__45641\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__10425\ : CascadeMux
    port map (
            O => \N__45638\,
            I => \N__45634\
        );

    \I__10424\ : InMux
    port map (
            O => \N__45637\,
            I => \N__45631\
        );

    \I__10423\ : InMux
    port map (
            O => \N__45634\,
            I => \N__45627\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__45631\,
            I => \N__45624\
        );

    \I__10421\ : InMux
    port map (
            O => \N__45630\,
            I => \N__45621\
        );

    \I__10420\ : LocalMux
    port map (
            O => \N__45627\,
            I => \N__45618\
        );

    \I__10419\ : Span4Mux_h
    port map (
            O => \N__45624\,
            I => \N__45615\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__45621\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__10417\ : Odrv12
    port map (
            O => \N__45618\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__10416\ : Odrv4
    port map (
            O => \N__45615\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__10415\ : InMux
    port map (
            O => \N__45608\,
            I => \N__45605\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__45605\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__10413\ : InMux
    port map (
            O => \N__45602\,
            I => \N__45599\
        );

    \I__10412\ : LocalMux
    port map (
            O => \N__45599\,
            I => \N__45596\
        );

    \I__10411\ : Odrv4
    port map (
            O => \N__45596\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__10410\ : InMux
    port map (
            O => \N__45593\,
            I => \N__45580\
        );

    \I__10409\ : InMux
    port map (
            O => \N__45592\,
            I => \N__45580\
        );

    \I__10408\ : InMux
    port map (
            O => \N__45591\,
            I => \N__45573\
        );

    \I__10407\ : InMux
    port map (
            O => \N__45590\,
            I => \N__45573\
        );

    \I__10406\ : InMux
    port map (
            O => \N__45589\,
            I => \N__45573\
        );

    \I__10405\ : InMux
    port map (
            O => \N__45588\,
            I => \N__45569\
        );

    \I__10404\ : InMux
    port map (
            O => \N__45587\,
            I => \N__45566\
        );

    \I__10403\ : InMux
    port map (
            O => \N__45586\,
            I => \N__45561\
        );

    \I__10402\ : InMux
    port map (
            O => \N__45585\,
            I => \N__45561\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__45580\,
            I => \N__45556\
        );

    \I__10400\ : LocalMux
    port map (
            O => \N__45573\,
            I => \N__45556\
        );

    \I__10399\ : InMux
    port map (
            O => \N__45572\,
            I => \N__45553\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__45569\,
            I => \N__45542\
        );

    \I__10397\ : LocalMux
    port map (
            O => \N__45566\,
            I => \N__45542\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__45561\,
            I => \N__45542\
        );

    \I__10395\ : Span4Mux_v
    port map (
            O => \N__45556\,
            I => \N__45537\
        );

    \I__10394\ : LocalMux
    port map (
            O => \N__45553\,
            I => \N__45537\
        );

    \I__10393\ : InMux
    port map (
            O => \N__45552\,
            I => \N__45528\
        );

    \I__10392\ : InMux
    port map (
            O => \N__45551\,
            I => \N__45528\
        );

    \I__10391\ : InMux
    port map (
            O => \N__45550\,
            I => \N__45528\
        );

    \I__10390\ : InMux
    port map (
            O => \N__45549\,
            I => \N__45528\
        );

    \I__10389\ : Span4Mux_v
    port map (
            O => \N__45542\,
            I => \N__45514\
        );

    \I__10388\ : Span4Mux_v
    port map (
            O => \N__45537\,
            I => \N__45509\
        );

    \I__10387\ : LocalMux
    port map (
            O => \N__45528\,
            I => \N__45509\
        );

    \I__10386\ : InMux
    port map (
            O => \N__45527\,
            I => \N__45492\
        );

    \I__10385\ : InMux
    port map (
            O => \N__45526\,
            I => \N__45492\
        );

    \I__10384\ : InMux
    port map (
            O => \N__45525\,
            I => \N__45492\
        );

    \I__10383\ : InMux
    port map (
            O => \N__45524\,
            I => \N__45492\
        );

    \I__10382\ : InMux
    port map (
            O => \N__45523\,
            I => \N__45492\
        );

    \I__10381\ : InMux
    port map (
            O => \N__45522\,
            I => \N__45492\
        );

    \I__10380\ : InMux
    port map (
            O => \N__45521\,
            I => \N__45492\
        );

    \I__10379\ : InMux
    port map (
            O => \N__45520\,
            I => \N__45492\
        );

    \I__10378\ : InMux
    port map (
            O => \N__45519\,
            I => \N__45489\
        );

    \I__10377\ : InMux
    port map (
            O => \N__45518\,
            I => \N__45484\
        );

    \I__10376\ : InMux
    port map (
            O => \N__45517\,
            I => \N__45484\
        );

    \I__10375\ : Odrv4
    port map (
            O => \N__45514\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10374\ : Odrv4
    port map (
            O => \N__45509\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10373\ : LocalMux
    port map (
            O => \N__45492\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__45489\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__45484\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10370\ : InMux
    port map (
            O => \N__45473\,
            I => \N__45469\
        );

    \I__10369\ : InMux
    port map (
            O => \N__45472\,
            I => \N__45466\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__45469\,
            I => \N__45462\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__45466\,
            I => \N__45459\
        );

    \I__10366\ : InMux
    port map (
            O => \N__45465\,
            I => \N__45456\
        );

    \I__10365\ : Span4Mux_h
    port map (
            O => \N__45462\,
            I => \N__45451\
        );

    \I__10364\ : Span4Mux_v
    port map (
            O => \N__45459\,
            I => \N__45451\
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__45456\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__10362\ : Odrv4
    port map (
            O => \N__45451\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__10361\ : CascadeMux
    port map (
            O => \N__45446\,
            I => \N__45443\
        );

    \I__10360\ : InMux
    port map (
            O => \N__45443\,
            I => \N__45440\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__45440\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__10358\ : InMux
    port map (
            O => \N__45437\,
            I => \N__45434\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__45434\,
            I => \N__45431\
        );

    \I__10356\ : Odrv4
    port map (
            O => \N__45431\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__10355\ : CascadeMux
    port map (
            O => \N__45428\,
            I => \N__45425\
        );

    \I__10354\ : InMux
    port map (
            O => \N__45425\,
            I => \N__45422\
        );

    \I__10353\ : LocalMux
    port map (
            O => \N__45422\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__10352\ : CascadeMux
    port map (
            O => \N__45419\,
            I => \N__45416\
        );

    \I__10351\ : InMux
    port map (
            O => \N__45416\,
            I => \N__45412\
        );

    \I__10350\ : CascadeMux
    port map (
            O => \N__45415\,
            I => \N__45409\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__45412\,
            I => \N__45405\
        );

    \I__10348\ : InMux
    port map (
            O => \N__45409\,
            I => \N__45402\
        );

    \I__10347\ : InMux
    port map (
            O => \N__45408\,
            I => \N__45399\
        );

    \I__10346\ : Span4Mux_h
    port map (
            O => \N__45405\,
            I => \N__45394\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__45402\,
            I => \N__45394\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__45399\,
            I => \N__45391\
        );

    \I__10343\ : Span4Mux_v
    port map (
            O => \N__45394\,
            I => \N__45388\
        );

    \I__10342\ : Odrv4
    port map (
            O => \N__45391\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__10341\ : Odrv4
    port map (
            O => \N__45388\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__10340\ : CascadeMux
    port map (
            O => \N__45383\,
            I => \N__45380\
        );

    \I__10339\ : InMux
    port map (
            O => \N__45380\,
            I => \N__45377\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__45377\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__10337\ : InMux
    port map (
            O => \N__45374\,
            I => \N__45371\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__45371\,
            I => \N__45368\
        );

    \I__10335\ : Span4Mux_h
    port map (
            O => \N__45368\,
            I => \N__45363\
        );

    \I__10334\ : InMux
    port map (
            O => \N__45367\,
            I => \N__45360\
        );

    \I__10333\ : InMux
    port map (
            O => \N__45366\,
            I => \N__45357\
        );

    \I__10332\ : Odrv4
    port map (
            O => \N__45363\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__45360\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__10330\ : LocalMux
    port map (
            O => \N__45357\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__10329\ : InMux
    port map (
            O => \N__45350\,
            I => \N__45347\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__45347\,
            I => \N__45344\
        );

    \I__10327\ : Odrv4
    port map (
            O => \N__45344\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\
        );

    \I__10326\ : CascadeMux
    port map (
            O => \N__45341\,
            I => \N__45338\
        );

    \I__10325\ : InMux
    port map (
            O => \N__45338\,
            I => \N__45335\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__45335\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__10323\ : CascadeMux
    port map (
            O => \N__45332\,
            I => \N__45328\
        );

    \I__10322\ : InMux
    port map (
            O => \N__45331\,
            I => \N__45322\
        );

    \I__10321\ : InMux
    port map (
            O => \N__45328\,
            I => \N__45322\
        );

    \I__10320\ : InMux
    port map (
            O => \N__45327\,
            I => \N__45319\
        );

    \I__10319\ : LocalMux
    port map (
            O => \N__45322\,
            I => \N__45316\
        );

    \I__10318\ : LocalMux
    port map (
            O => \N__45319\,
            I => \N__45313\
        );

    \I__10317\ : Span4Mux_h
    port map (
            O => \N__45316\,
            I => \N__45310\
        );

    \I__10316\ : Span4Mux_h
    port map (
            O => \N__45313\,
            I => \N__45307\
        );

    \I__10315\ : Odrv4
    port map (
            O => \N__45310\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__10314\ : Odrv4
    port map (
            O => \N__45307\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__10313\ : CascadeMux
    port map (
            O => \N__45302\,
            I => \N__45299\
        );

    \I__10312\ : InMux
    port map (
            O => \N__45299\,
            I => \N__45296\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__45296\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__10310\ : CascadeMux
    port map (
            O => \N__45293\,
            I => \N__45290\
        );

    \I__10309\ : InMux
    port map (
            O => \N__45290\,
            I => \N__45287\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__45287\,
            I => \N__45282\
        );

    \I__10307\ : InMux
    port map (
            O => \N__45286\,
            I => \N__45279\
        );

    \I__10306\ : InMux
    port map (
            O => \N__45285\,
            I => \N__45276\
        );

    \I__10305\ : Span4Mux_h
    port map (
            O => \N__45282\,
            I => \N__45271\
        );

    \I__10304\ : LocalMux
    port map (
            O => \N__45279\,
            I => \N__45271\
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__45276\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__10302\ : Odrv4
    port map (
            O => \N__45271\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__10301\ : InMux
    port map (
            O => \N__45266\,
            I => \N__45263\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__45263\,
            I => \N__45260\
        );

    \I__10299\ : Odrv4
    port map (
            O => \N__45260\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__10298\ : CascadeMux
    port map (
            O => \N__45257\,
            I => \N__45254\
        );

    \I__10297\ : InMux
    port map (
            O => \N__45254\,
            I => \N__45251\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__45251\,
            I => \N__45246\
        );

    \I__10295\ : InMux
    port map (
            O => \N__45250\,
            I => \N__45243\
        );

    \I__10294\ : InMux
    port map (
            O => \N__45249\,
            I => \N__45240\
        );

    \I__10293\ : Span4Mux_v
    port map (
            O => \N__45246\,
            I => \N__45235\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__45243\,
            I => \N__45235\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__45240\,
            I => \N__45232\
        );

    \I__10290\ : Span4Mux_h
    port map (
            O => \N__45235\,
            I => \N__45229\
        );

    \I__10289\ : Odrv4
    port map (
            O => \N__45232\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__10288\ : Odrv4
    port map (
            O => \N__45229\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__10287\ : CascadeMux
    port map (
            O => \N__45224\,
            I => \N__45221\
        );

    \I__10286\ : InMux
    port map (
            O => \N__45221\,
            I => \N__45218\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__45218\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__10284\ : CascadeMux
    port map (
            O => \N__45215\,
            I => \N__45212\
        );

    \I__10283\ : InMux
    port map (
            O => \N__45212\,
            I => \N__45207\
        );

    \I__10282\ : InMux
    port map (
            O => \N__45211\,
            I => \N__45204\
        );

    \I__10281\ : InMux
    port map (
            O => \N__45210\,
            I => \N__45201\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__45207\,
            I => \N__45198\
        );

    \I__10279\ : LocalMux
    port map (
            O => \N__45204\,
            I => \N__45195\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__45201\,
            I => \N__45192\
        );

    \I__10277\ : Span4Mux_v
    port map (
            O => \N__45198\,
            I => \N__45187\
        );

    \I__10276\ : Span4Mux_h
    port map (
            O => \N__45195\,
            I => \N__45187\
        );

    \I__10275\ : Span4Mux_h
    port map (
            O => \N__45192\,
            I => \N__45184\
        );

    \I__10274\ : Odrv4
    port map (
            O => \N__45187\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__10273\ : Odrv4
    port map (
            O => \N__45184\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__10272\ : InMux
    port map (
            O => \N__45179\,
            I => \N__45176\
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__45176\,
            I => \N__45173\
        );

    \I__10270\ : Odrv12
    port map (
            O => \N__45173\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\
        );

    \I__10269\ : InMux
    port map (
            O => \N__45170\,
            I => \N__45165\
        );

    \I__10268\ : InMux
    port map (
            O => \N__45169\,
            I => \N__45162\
        );

    \I__10267\ : InMux
    port map (
            O => \N__45168\,
            I => \N__45159\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__45165\,
            I => \N__45156\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__45162\,
            I => \N__45153\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__45159\,
            I => \N__45150\
        );

    \I__10263\ : Sp12to4
    port map (
            O => \N__45156\,
            I => \N__45147\
        );

    \I__10262\ : Span4Mux_v
    port map (
            O => \N__45153\,
            I => \N__45144\
        );

    \I__10261\ : Span4Mux_h
    port map (
            O => \N__45150\,
            I => \N__45141\
        );

    \I__10260\ : Odrv12
    port map (
            O => \N__45147\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10259\ : Odrv4
    port map (
            O => \N__45144\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10258\ : Odrv4
    port map (
            O => \N__45141\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10257\ : InMux
    port map (
            O => \N__45134\,
            I => \N__45131\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__45131\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__10255\ : InMux
    port map (
            O => \N__45128\,
            I => \N__45122\
        );

    \I__10254\ : InMux
    port map (
            O => \N__45127\,
            I => \N__45122\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__45122\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\
        );

    \I__10252\ : CEMux
    port map (
            O => \N__45119\,
            I => \N__45092\
        );

    \I__10251\ : CEMux
    port map (
            O => \N__45118\,
            I => \N__45092\
        );

    \I__10250\ : CEMux
    port map (
            O => \N__45117\,
            I => \N__45092\
        );

    \I__10249\ : CEMux
    port map (
            O => \N__45116\,
            I => \N__45092\
        );

    \I__10248\ : CEMux
    port map (
            O => \N__45115\,
            I => \N__45092\
        );

    \I__10247\ : CEMux
    port map (
            O => \N__45114\,
            I => \N__45092\
        );

    \I__10246\ : CEMux
    port map (
            O => \N__45113\,
            I => \N__45092\
        );

    \I__10245\ : CEMux
    port map (
            O => \N__45112\,
            I => \N__45092\
        );

    \I__10244\ : CEMux
    port map (
            O => \N__45111\,
            I => \N__45092\
        );

    \I__10243\ : GlobalMux
    port map (
            O => \N__45092\,
            I => \N__45089\
        );

    \I__10242\ : gio2CtrlBuf
    port map (
            O => \N__45089\,
            I => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \I__10241\ : InMux
    port map (
            O => \N__45086\,
            I => \N__45082\
        );

    \I__10240\ : CascadeMux
    port map (
            O => \N__45085\,
            I => \N__45078\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__45082\,
            I => \N__45075\
        );

    \I__10238\ : InMux
    port map (
            O => \N__45081\,
            I => \N__45072\
        );

    \I__10237\ : InMux
    port map (
            O => \N__45078\,
            I => \N__45069\
        );

    \I__10236\ : Span4Mux_h
    port map (
            O => \N__45075\,
            I => \N__45062\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__45072\,
            I => \N__45062\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__45069\,
            I => \N__45062\
        );

    \I__10233\ : Odrv4
    port map (
            O => \N__45062\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__10232\ : CascadeMux
    port map (
            O => \N__45059\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__10231\ : InMux
    port map (
            O => \N__45056\,
            I => \N__45052\
        );

    \I__10230\ : CascadeMux
    port map (
            O => \N__45055\,
            I => \N__45049\
        );

    \I__10229\ : LocalMux
    port map (
            O => \N__45052\,
            I => \N__45046\
        );

    \I__10228\ : InMux
    port map (
            O => \N__45049\,
            I => \N__45043\
        );

    \I__10227\ : Span4Mux_v
    port map (
            O => \N__45046\,
            I => \N__45038\
        );

    \I__10226\ : LocalMux
    port map (
            O => \N__45043\,
            I => \N__45038\
        );

    \I__10225\ : Odrv4
    port map (
            O => \N__45038\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__10224\ : InMux
    port map (
            O => \N__45035\,
            I => \N__45032\
        );

    \I__10223\ : LocalMux
    port map (
            O => \N__45032\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__10222\ : InMux
    port map (
            O => \N__45029\,
            I => \N__45025\
        );

    \I__10221\ : CascadeMux
    port map (
            O => \N__45028\,
            I => \N__45020\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__45025\,
            I => \N__45017\
        );

    \I__10219\ : InMux
    port map (
            O => \N__45024\,
            I => \N__45012\
        );

    \I__10218\ : InMux
    port map (
            O => \N__45023\,
            I => \N__45012\
        );

    \I__10217\ : InMux
    port map (
            O => \N__45020\,
            I => \N__45009\
        );

    \I__10216\ : Span4Mux_v
    port map (
            O => \N__45017\,
            I => \N__45004\
        );

    \I__10215\ : LocalMux
    port map (
            O => \N__45012\,
            I => \N__45004\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__45009\,
            I => \N__44998\
        );

    \I__10213\ : Span4Mux_v
    port map (
            O => \N__45004\,
            I => \N__44998\
        );

    \I__10212\ : InMux
    port map (
            O => \N__45003\,
            I => \N__44995\
        );

    \I__10211\ : Odrv4
    port map (
            O => \N__44998\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__44995\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__10209\ : CascadeMux
    port map (
            O => \N__44990\,
            I => \N__44982\
        );

    \I__10208\ : CascadeMux
    port map (
            O => \N__44989\,
            I => \N__44978\
        );

    \I__10207\ : CascadeMux
    port map (
            O => \N__44988\,
            I => \N__44974\
        );

    \I__10206\ : InMux
    port map (
            O => \N__44987\,
            I => \N__44953\
        );

    \I__10205\ : InMux
    port map (
            O => \N__44986\,
            I => \N__44953\
        );

    \I__10204\ : InMux
    port map (
            O => \N__44985\,
            I => \N__44938\
        );

    \I__10203\ : InMux
    port map (
            O => \N__44982\,
            I => \N__44938\
        );

    \I__10202\ : InMux
    port map (
            O => \N__44981\,
            I => \N__44938\
        );

    \I__10201\ : InMux
    port map (
            O => \N__44978\,
            I => \N__44938\
        );

    \I__10200\ : InMux
    port map (
            O => \N__44977\,
            I => \N__44938\
        );

    \I__10199\ : InMux
    port map (
            O => \N__44974\,
            I => \N__44938\
        );

    \I__10198\ : InMux
    port map (
            O => \N__44973\,
            I => \N__44938\
        );

    \I__10197\ : CascadeMux
    port map (
            O => \N__44972\,
            I => \N__44931\
        );

    \I__10196\ : CascadeMux
    port map (
            O => \N__44971\,
            I => \N__44927\
        );

    \I__10195\ : CascadeMux
    port map (
            O => \N__44970\,
            I => \N__44923\
        );

    \I__10194\ : CascadeMux
    port map (
            O => \N__44969\,
            I => \N__44919\
        );

    \I__10193\ : CascadeMux
    port map (
            O => \N__44968\,
            I => \N__44914\
        );

    \I__10192\ : CascadeMux
    port map (
            O => \N__44967\,
            I => \N__44910\
        );

    \I__10191\ : CascadeMux
    port map (
            O => \N__44966\,
            I => \N__44906\
        );

    \I__10190\ : InMux
    port map (
            O => \N__44965\,
            I => \N__44902\
        );

    \I__10189\ : InMux
    port map (
            O => \N__44964\,
            I => \N__44895\
        );

    \I__10188\ : InMux
    port map (
            O => \N__44963\,
            I => \N__44895\
        );

    \I__10187\ : InMux
    port map (
            O => \N__44962\,
            I => \N__44895\
        );

    \I__10186\ : InMux
    port map (
            O => \N__44961\,
            I => \N__44882\
        );

    \I__10185\ : InMux
    port map (
            O => \N__44960\,
            I => \N__44882\
        );

    \I__10184\ : InMux
    port map (
            O => \N__44959\,
            I => \N__44882\
        );

    \I__10183\ : InMux
    port map (
            O => \N__44958\,
            I => \N__44882\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__44953\,
            I => \N__44877\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__44938\,
            I => \N__44877\
        );

    \I__10180\ : InMux
    port map (
            O => \N__44937\,
            I => \N__44868\
        );

    \I__10179\ : InMux
    port map (
            O => \N__44936\,
            I => \N__44868\
        );

    \I__10178\ : InMux
    port map (
            O => \N__44935\,
            I => \N__44868\
        );

    \I__10177\ : InMux
    port map (
            O => \N__44934\,
            I => \N__44868\
        );

    \I__10176\ : InMux
    port map (
            O => \N__44931\,
            I => \N__44851\
        );

    \I__10175\ : InMux
    port map (
            O => \N__44930\,
            I => \N__44851\
        );

    \I__10174\ : InMux
    port map (
            O => \N__44927\,
            I => \N__44851\
        );

    \I__10173\ : InMux
    port map (
            O => \N__44926\,
            I => \N__44851\
        );

    \I__10172\ : InMux
    port map (
            O => \N__44923\,
            I => \N__44851\
        );

    \I__10171\ : InMux
    port map (
            O => \N__44922\,
            I => \N__44851\
        );

    \I__10170\ : InMux
    port map (
            O => \N__44919\,
            I => \N__44851\
        );

    \I__10169\ : InMux
    port map (
            O => \N__44918\,
            I => \N__44851\
        );

    \I__10168\ : InMux
    port map (
            O => \N__44917\,
            I => \N__44836\
        );

    \I__10167\ : InMux
    port map (
            O => \N__44914\,
            I => \N__44836\
        );

    \I__10166\ : InMux
    port map (
            O => \N__44913\,
            I => \N__44836\
        );

    \I__10165\ : InMux
    port map (
            O => \N__44910\,
            I => \N__44836\
        );

    \I__10164\ : InMux
    port map (
            O => \N__44909\,
            I => \N__44836\
        );

    \I__10163\ : InMux
    port map (
            O => \N__44906\,
            I => \N__44836\
        );

    \I__10162\ : InMux
    port map (
            O => \N__44905\,
            I => \N__44836\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__44902\,
            I => \N__44826\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__44895\,
            I => \N__44826\
        );

    \I__10159\ : InMux
    port map (
            O => \N__44894\,
            I => \N__44817\
        );

    \I__10158\ : InMux
    port map (
            O => \N__44893\,
            I => \N__44817\
        );

    \I__10157\ : InMux
    port map (
            O => \N__44892\,
            I => \N__44817\
        );

    \I__10156\ : InMux
    port map (
            O => \N__44891\,
            I => \N__44817\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__44882\,
            I => \N__44810\
        );

    \I__10154\ : Span4Mux_v
    port map (
            O => \N__44877\,
            I => \N__44801\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__44868\,
            I => \N__44801\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__44851\,
            I => \N__44801\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__44836\,
            I => \N__44801\
        );

    \I__10150\ : InMux
    port map (
            O => \N__44835\,
            I => \N__44798\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44834\,
            I => \N__44793\
        );

    \I__10148\ : InMux
    port map (
            O => \N__44833\,
            I => \N__44793\
        );

    \I__10147\ : InMux
    port map (
            O => \N__44832\,
            I => \N__44790\
        );

    \I__10146\ : InMux
    port map (
            O => \N__44831\,
            I => \N__44787\
        );

    \I__10145\ : Span4Mux_v
    port map (
            O => \N__44826\,
            I => \N__44782\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__44817\,
            I => \N__44779\
        );

    \I__10143\ : InMux
    port map (
            O => \N__44816\,
            I => \N__44776\
        );

    \I__10142\ : InMux
    port map (
            O => \N__44815\,
            I => \N__44771\
        );

    \I__10141\ : InMux
    port map (
            O => \N__44814\,
            I => \N__44771\
        );

    \I__10140\ : InMux
    port map (
            O => \N__44813\,
            I => \N__44768\
        );

    \I__10139\ : Span4Mux_v
    port map (
            O => \N__44810\,
            I => \N__44763\
        );

    \I__10138\ : Span4Mux_v
    port map (
            O => \N__44801\,
            I => \N__44763\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__44798\,
            I => \N__44754\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__44793\,
            I => \N__44754\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__44790\,
            I => \N__44754\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__44787\,
            I => \N__44754\
        );

    \I__10133\ : InMux
    port map (
            O => \N__44786\,
            I => \N__44751\
        );

    \I__10132\ : InMux
    port map (
            O => \N__44785\,
            I => \N__44748\
        );

    \I__10131\ : Span4Mux_h
    port map (
            O => \N__44782\,
            I => \N__44735\
        );

    \I__10130\ : Span4Mux_v
    port map (
            O => \N__44779\,
            I => \N__44735\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__44776\,
            I => \N__44735\
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__44771\,
            I => \N__44735\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__44768\,
            I => \N__44735\
        );

    \I__10126\ : Sp12to4
    port map (
            O => \N__44763\,
            I => \N__44730\
        );

    \I__10125\ : Span12Mux_s11_v
    port map (
            O => \N__44754\,
            I => \N__44730\
        );

    \I__10124\ : LocalMux
    port map (
            O => \N__44751\,
            I => \N__44727\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__44748\,
            I => \N__44724\
        );

    \I__10122\ : InMux
    port map (
            O => \N__44747\,
            I => \N__44721\
        );

    \I__10121\ : CascadeMux
    port map (
            O => \N__44746\,
            I => \N__44717\
        );

    \I__10120\ : Sp12to4
    port map (
            O => \N__44735\,
            I => \N__44705\
        );

    \I__10119\ : Span12Mux_h
    port map (
            O => \N__44730\,
            I => \N__44702\
        );

    \I__10118\ : Span4Mux_s1_h
    port map (
            O => \N__44727\,
            I => \N__44695\
        );

    \I__10117\ : Span4Mux_s1_v
    port map (
            O => \N__44724\,
            I => \N__44695\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__44721\,
            I => \N__44695\
        );

    \I__10115\ : InMux
    port map (
            O => \N__44720\,
            I => \N__44688\
        );

    \I__10114\ : InMux
    port map (
            O => \N__44717\,
            I => \N__44688\
        );

    \I__10113\ : InMux
    port map (
            O => \N__44716\,
            I => \N__44688\
        );

    \I__10112\ : InMux
    port map (
            O => \N__44715\,
            I => \N__44685\
        );

    \I__10111\ : InMux
    port map (
            O => \N__44714\,
            I => \N__44678\
        );

    \I__10110\ : InMux
    port map (
            O => \N__44713\,
            I => \N__44678\
        );

    \I__10109\ : InMux
    port map (
            O => \N__44712\,
            I => \N__44678\
        );

    \I__10108\ : InMux
    port map (
            O => \N__44711\,
            I => \N__44669\
        );

    \I__10107\ : InMux
    port map (
            O => \N__44710\,
            I => \N__44669\
        );

    \I__10106\ : InMux
    port map (
            O => \N__44709\,
            I => \N__44669\
        );

    \I__10105\ : InMux
    port map (
            O => \N__44708\,
            I => \N__44669\
        );

    \I__10104\ : Span12Mux_v
    port map (
            O => \N__44705\,
            I => \N__44660\
        );

    \I__10103\ : Span12Mux_h
    port map (
            O => \N__44702\,
            I => \N__44660\
        );

    \I__10102\ : Sp12to4
    port map (
            O => \N__44695\,
            I => \N__44660\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__44688\,
            I => \N__44660\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__44685\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__44678\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__44669\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10097\ : Odrv12
    port map (
            O => \N__44660\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10096\ : CascadeMux
    port map (
            O => \N__44651\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\
        );

    \I__10095\ : CascadeMux
    port map (
            O => \N__44648\,
            I => \N__44645\
        );

    \I__10094\ : InMux
    port map (
            O => \N__44645\,
            I => \N__44642\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__44642\,
            I => \N__44638\
        );

    \I__10092\ : InMux
    port map (
            O => \N__44641\,
            I => \N__44635\
        );

    \I__10091\ : Span4Mux_h
    port map (
            O => \N__44638\,
            I => \N__44632\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__44635\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__10089\ : Odrv4
    port map (
            O => \N__44632\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__10088\ : InMux
    port map (
            O => \N__44627\,
            I => \N__44624\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__44624\,
            I => \N__44620\
        );

    \I__10086\ : InMux
    port map (
            O => \N__44623\,
            I => \N__44617\
        );

    \I__10085\ : Span4Mux_v
    port map (
            O => \N__44620\,
            I => \N__44612\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__44617\,
            I => \N__44612\
        );

    \I__10083\ : Span4Mux_h
    port map (
            O => \N__44612\,
            I => \N__44609\
        );

    \I__10082\ : Odrv4
    port map (
            O => \N__44609\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__10081\ : InMux
    port map (
            O => \N__44606\,
            I => \N__44602\
        );

    \I__10080\ : InMux
    port map (
            O => \N__44605\,
            I => \N__44599\
        );

    \I__10079\ : LocalMux
    port map (
            O => \N__44602\,
            I => \N__44595\
        );

    \I__10078\ : LocalMux
    port map (
            O => \N__44599\,
            I => \N__44592\
        );

    \I__10077\ : InMux
    port map (
            O => \N__44598\,
            I => \N__44589\
        );

    \I__10076\ : Span4Mux_h
    port map (
            O => \N__44595\,
            I => \N__44586\
        );

    \I__10075\ : Odrv12
    port map (
            O => \N__44592\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__44589\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10073\ : Odrv4
    port map (
            O => \N__44586\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10072\ : CascadeMux
    port map (
            O => \N__44579\,
            I => \N__44576\
        );

    \I__10071\ : InMux
    port map (
            O => \N__44576\,
            I => \N__44573\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__44573\,
            I => \N__44570\
        );

    \I__10069\ : Span4Mux_h
    port map (
            O => \N__44570\,
            I => \N__44567\
        );

    \I__10068\ : Odrv4
    port map (
            O => \N__44567\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__10067\ : InMux
    port map (
            O => \N__44564\,
            I => \N__44561\
        );

    \I__10066\ : LocalMux
    port map (
            O => \N__44561\,
            I => \N__44558\
        );

    \I__10065\ : Span4Mux_v
    port map (
            O => \N__44558\,
            I => \N__44555\
        );

    \I__10064\ : Odrv4
    port map (
            O => \N__44555\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__10063\ : InMux
    port map (
            O => \N__44552\,
            I => \N__44548\
        );

    \I__10062\ : InMux
    port map (
            O => \N__44551\,
            I => \N__44545\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__44548\,
            I => \N__44542\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__44545\,
            I => \N__44538\
        );

    \I__10059\ : Span4Mux_h
    port map (
            O => \N__44542\,
            I => \N__44535\
        );

    \I__10058\ : InMux
    port map (
            O => \N__44541\,
            I => \N__44532\
        );

    \I__10057\ : Odrv12
    port map (
            O => \N__44538\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__10056\ : Odrv4
    port map (
            O => \N__44535\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__10055\ : LocalMux
    port map (
            O => \N__44532\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__10054\ : InMux
    port map (
            O => \N__44525\,
            I => \N__44522\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__44522\,
            I => \N__44519\
        );

    \I__10052\ : Odrv12
    port map (
            O => \N__44519\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\
        );

    \I__10051\ : InMux
    port map (
            O => \N__44516\,
            I => \N__44513\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__44513\,
            I => \N__44509\
        );

    \I__10049\ : InMux
    port map (
            O => \N__44512\,
            I => \N__44506\
        );

    \I__10048\ : Span4Mux_v
    port map (
            O => \N__44509\,
            I => \N__44500\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__44506\,
            I => \N__44500\
        );

    \I__10046\ : InMux
    port map (
            O => \N__44505\,
            I => \N__44496\
        );

    \I__10045\ : Span4Mux_v
    port map (
            O => \N__44500\,
            I => \N__44493\
        );

    \I__10044\ : InMux
    port map (
            O => \N__44499\,
            I => \N__44490\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__44496\,
            I => \N__44487\
        );

    \I__10042\ : Odrv4
    port map (
            O => \N__44493\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__44490\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__10040\ : Odrv4
    port map (
            O => \N__44487\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__10039\ : InMux
    port map (
            O => \N__44480\,
            I => \N__44477\
        );

    \I__10038\ : LocalMux
    port map (
            O => \N__44477\,
            I => \N__44474\
        );

    \I__10037\ : Span4Mux_v
    port map (
            O => \N__44474\,
            I => \N__44470\
        );

    \I__10036\ : InMux
    port map (
            O => \N__44473\,
            I => \N__44467\
        );

    \I__10035\ : Span4Mux_v
    port map (
            O => \N__44470\,
            I => \N__44461\
        );

    \I__10034\ : LocalMux
    port map (
            O => \N__44467\,
            I => \N__44461\
        );

    \I__10033\ : InMux
    port map (
            O => \N__44466\,
            I => \N__44458\
        );

    \I__10032\ : Span4Mux_h
    port map (
            O => \N__44461\,
            I => \N__44455\
        );

    \I__10031\ : LocalMux
    port map (
            O => \N__44458\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10030\ : Odrv4
    port map (
            O => \N__44455\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10029\ : CascadeMux
    port map (
            O => \N__44450\,
            I => \N__44447\
        );

    \I__10028\ : InMux
    port map (
            O => \N__44447\,
            I => \N__44444\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__44444\,
            I => \N__44441\
        );

    \I__10026\ : Odrv12
    port map (
            O => \N__44441\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt24\
        );

    \I__10025\ : InMux
    port map (
            O => \N__44438\,
            I => \N__44431\
        );

    \I__10024\ : InMux
    port map (
            O => \N__44437\,
            I => \N__44431\
        );

    \I__10023\ : InMux
    port map (
            O => \N__44436\,
            I => \N__44428\
        );

    \I__10022\ : LocalMux
    port map (
            O => \N__44431\,
            I => \N__44425\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__44428\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__10020\ : Odrv12
    port map (
            O => \N__44425\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__10019\ : CascadeMux
    port map (
            O => \N__44420\,
            I => \N__44417\
        );

    \I__10018\ : InMux
    port map (
            O => \N__44417\,
            I => \N__44411\
        );

    \I__10017\ : InMux
    port map (
            O => \N__44416\,
            I => \N__44411\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__44411\,
            I => \N__44407\
        );

    \I__10015\ : InMux
    port map (
            O => \N__44410\,
            I => \N__44404\
        );

    \I__10014\ : Span4Mux_v
    port map (
            O => \N__44407\,
            I => \N__44401\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__44404\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__10012\ : Odrv4
    port map (
            O => \N__44401\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__10011\ : InMux
    port map (
            O => \N__44396\,
            I => \N__44393\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__44393\,
            I => \N__44390\
        );

    \I__10009\ : Odrv12
    port map (
            O => \N__44390\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\
        );

    \I__10008\ : InMux
    port map (
            O => \N__44387\,
            I => \N__44382\
        );

    \I__10007\ : InMux
    port map (
            O => \N__44386\,
            I => \N__44379\
        );

    \I__10006\ : InMux
    port map (
            O => \N__44385\,
            I => \N__44376\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__44382\,
            I => \N__44371\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__44379\,
            I => \N__44371\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__44376\,
            I => \N__44368\
        );

    \I__10002\ : Span4Mux_v
    port map (
            O => \N__44371\,
            I => \N__44365\
        );

    \I__10001\ : Span4Mux_v
    port map (
            O => \N__44368\,
            I => \N__44359\
        );

    \I__10000\ : Span4Mux_h
    port map (
            O => \N__44365\,
            I => \N__44359\
        );

    \I__9999\ : InMux
    port map (
            O => \N__44364\,
            I => \N__44356\
        );

    \I__9998\ : Odrv4
    port map (
            O => \N__44359\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__9997\ : LocalMux
    port map (
            O => \N__44356\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__9996\ : InMux
    port map (
            O => \N__44351\,
            I => \N__44348\
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__44348\,
            I => \N__44345\
        );

    \I__9994\ : Span4Mux_v
    port map (
            O => \N__44345\,
            I => \N__44342\
        );

    \I__9993\ : Span4Mux_h
    port map (
            O => \N__44342\,
            I => \N__44337\
        );

    \I__9992\ : InMux
    port map (
            O => \N__44341\,
            I => \N__44334\
        );

    \I__9991\ : InMux
    port map (
            O => \N__44340\,
            I => \N__44331\
        );

    \I__9990\ : Span4Mux_h
    port map (
            O => \N__44337\,
            I => \N__44328\
        );

    \I__9989\ : LocalMux
    port map (
            O => \N__44334\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__44331\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__9987\ : Odrv4
    port map (
            O => \N__44328\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__9986\ : InMux
    port map (
            O => \N__44321\,
            I => \N__44315\
        );

    \I__9985\ : InMux
    port map (
            O => \N__44320\,
            I => \N__44315\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__44315\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\
        );

    \I__9983\ : InMux
    port map (
            O => \N__44312\,
            I => \N__44309\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__44309\,
            I => \N__44306\
        );

    \I__9981\ : Span4Mux_h
    port map (
            O => \N__44306\,
            I => \N__44302\
        );

    \I__9980\ : InMux
    port map (
            O => \N__44305\,
            I => \N__44299\
        );

    \I__9979\ : Span4Mux_v
    port map (
            O => \N__44302\,
            I => \N__44295\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__44299\,
            I => \N__44292\
        );

    \I__9977\ : InMux
    port map (
            O => \N__44298\,
            I => \N__44289\
        );

    \I__9976\ : Span4Mux_h
    port map (
            O => \N__44295\,
            I => \N__44286\
        );

    \I__9975\ : Span4Mux_s2_v
    port map (
            O => \N__44292\,
            I => \N__44283\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__44289\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__9973\ : Odrv4
    port map (
            O => \N__44286\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__9972\ : Odrv4
    port map (
            O => \N__44283\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__9971\ : InMux
    port map (
            O => \N__44276\,
            I => \N__44273\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__44273\,
            I => \N__44268\
        );

    \I__9969\ : InMux
    port map (
            O => \N__44272\,
            I => \N__44265\
        );

    \I__9968\ : InMux
    port map (
            O => \N__44271\,
            I => \N__44262\
        );

    \I__9967\ : Span4Mux_v
    port map (
            O => \N__44268\,
            I => \N__44257\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__44265\,
            I => \N__44257\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__44262\,
            I => \N__44253\
        );

    \I__9964\ : Span4Mux_v
    port map (
            O => \N__44257\,
            I => \N__44250\
        );

    \I__9963\ : CascadeMux
    port map (
            O => \N__44256\,
            I => \N__44247\
        );

    \I__9962\ : Span4Mux_v
    port map (
            O => \N__44253\,
            I => \N__44244\
        );

    \I__9961\ : Span4Mux_h
    port map (
            O => \N__44250\,
            I => \N__44241\
        );

    \I__9960\ : InMux
    port map (
            O => \N__44247\,
            I => \N__44238\
        );

    \I__9959\ : Odrv4
    port map (
            O => \N__44244\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__9958\ : Odrv4
    port map (
            O => \N__44241\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__44238\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__9956\ : CascadeMux
    port map (
            O => \N__44231\,
            I => \N__44228\
        );

    \I__9955\ : InMux
    port map (
            O => \N__44228\,
            I => \N__44222\
        );

    \I__9954\ : InMux
    port map (
            O => \N__44227\,
            I => \N__44222\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__44222\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\
        );

    \I__9952\ : InMux
    port map (
            O => \N__44219\,
            I => \N__44216\
        );

    \I__9951\ : LocalMux
    port map (
            O => \N__44216\,
            I => \N__44213\
        );

    \I__9950\ : Odrv4
    port map (
            O => \N__44213\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\
        );

    \I__9949\ : InMux
    port map (
            O => \N__44210\,
            I => \N__44204\
        );

    \I__9948\ : InMux
    port map (
            O => \N__44209\,
            I => \N__44204\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__44204\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\
        );

    \I__9946\ : CascadeMux
    port map (
            O => \N__44201\,
            I => \N__44197\
        );

    \I__9945\ : InMux
    port map (
            O => \N__44200\,
            I => \N__44192\
        );

    \I__9944\ : InMux
    port map (
            O => \N__44197\,
            I => \N__44192\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__44192\,
            I => \N__44188\
        );

    \I__9942\ : InMux
    port map (
            O => \N__44191\,
            I => \N__44185\
        );

    \I__9941\ : Span4Mux_v
    port map (
            O => \N__44188\,
            I => \N__44182\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__44185\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__9939\ : Odrv4
    port map (
            O => \N__44182\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__9938\ : CascadeMux
    port map (
            O => \N__44177\,
            I => \N__44173\
        );

    \I__9937\ : InMux
    port map (
            O => \N__44176\,
            I => \N__44168\
        );

    \I__9936\ : InMux
    port map (
            O => \N__44173\,
            I => \N__44168\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__44168\,
            I => \N__44164\
        );

    \I__9934\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44161\
        );

    \I__9933\ : Span4Mux_h
    port map (
            O => \N__44164\,
            I => \N__44158\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__44161\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__9931\ : Odrv4
    port map (
            O => \N__44158\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__9930\ : CascadeMux
    port map (
            O => \N__44153\,
            I => \N__44150\
        );

    \I__9929\ : InMux
    port map (
            O => \N__44150\,
            I => \N__44147\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__44147\,
            I => \N__44144\
        );

    \I__9927\ : Odrv12
    port map (
            O => \N__44144\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__9926\ : InMux
    port map (
            O => \N__44141\,
            I => \N__44133\
        );

    \I__9925\ : InMux
    port map (
            O => \N__44140\,
            I => \N__44133\
        );

    \I__9924\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44130\
        );

    \I__9923\ : InMux
    port map (
            O => \N__44138\,
            I => \N__44127\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__44133\,
            I => \N__44122\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__44130\,
            I => \N__44122\
        );

    \I__9920\ : LocalMux
    port map (
            O => \N__44127\,
            I => \N__44119\
        );

    \I__9919\ : Span4Mux_v
    port map (
            O => \N__44122\,
            I => \N__44116\
        );

    \I__9918\ : Odrv12
    port map (
            O => \N__44119\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__9917\ : Odrv4
    port map (
            O => \N__44116\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__9916\ : InMux
    port map (
            O => \N__44111\,
            I => \N__44108\
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__44108\,
            I => \N__44105\
        );

    \I__9914\ : Span4Mux_v
    port map (
            O => \N__44105\,
            I => \N__44102\
        );

    \I__9913\ : Span4Mux_v
    port map (
            O => \N__44102\,
            I => \N__44098\
        );

    \I__9912\ : InMux
    port map (
            O => \N__44101\,
            I => \N__44095\
        );

    \I__9911\ : Odrv4
    port map (
            O => \N__44098\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__44095\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__9909\ : CascadeMux
    port map (
            O => \N__44090\,
            I => \N__44087\
        );

    \I__9908\ : InMux
    port map (
            O => \N__44087\,
            I => \N__44083\
        );

    \I__9907\ : InMux
    port map (
            O => \N__44086\,
            I => \N__44080\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__44083\,
            I => \N__44074\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__44080\,
            I => \N__44074\
        );

    \I__9904\ : InMux
    port map (
            O => \N__44079\,
            I => \N__44071\
        );

    \I__9903\ : Span4Mux_h
    port map (
            O => \N__44074\,
            I => \N__44068\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__44071\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__9901\ : Odrv4
    port map (
            O => \N__44068\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__9900\ : InMux
    port map (
            O => \N__44063\,
            I => \N__44060\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__44060\,
            I => \N__44055\
        );

    \I__9898\ : InMux
    port map (
            O => \N__44059\,
            I => \N__44052\
        );

    \I__9897\ : InMux
    port map (
            O => \N__44058\,
            I => \N__44049\
        );

    \I__9896\ : Span4Mux_v
    port map (
            O => \N__44055\,
            I => \N__44044\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__44052\,
            I => \N__44044\
        );

    \I__9894\ : LocalMux
    port map (
            O => \N__44049\,
            I => \N__44041\
        );

    \I__9893\ : Span4Mux_h
    port map (
            O => \N__44044\,
            I => \N__44038\
        );

    \I__9892\ : Span4Mux_h
    port map (
            O => \N__44041\,
            I => \N__44034\
        );

    \I__9891\ : Span4Mux_v
    port map (
            O => \N__44038\,
            I => \N__44031\
        );

    \I__9890\ : InMux
    port map (
            O => \N__44037\,
            I => \N__44028\
        );

    \I__9889\ : Odrv4
    port map (
            O => \N__44034\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__9888\ : Odrv4
    port map (
            O => \N__44031\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__44028\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__9886\ : InMux
    port map (
            O => \N__44021\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__9885\ : CascadeMux
    port map (
            O => \N__44018\,
            I => \N__44015\
        );

    \I__9884\ : InMux
    port map (
            O => \N__44015\,
            I => \N__44011\
        );

    \I__9883\ : InMux
    port map (
            O => \N__44014\,
            I => \N__44008\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__44011\,
            I => \N__44004\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__44008\,
            I => \N__44001\
        );

    \I__9880\ : InMux
    port map (
            O => \N__44007\,
            I => \N__43998\
        );

    \I__9879\ : Span4Mux_h
    port map (
            O => \N__44004\,
            I => \N__43995\
        );

    \I__9878\ : Span4Mux_h
    port map (
            O => \N__44001\,
            I => \N__43992\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__43998\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__9876\ : Odrv4
    port map (
            O => \N__43995\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__9875\ : Odrv4
    port map (
            O => \N__43992\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__9874\ : InMux
    port map (
            O => \N__43985\,
            I => \N__43980\
        );

    \I__9873\ : InMux
    port map (
            O => \N__43984\,
            I => \N__43977\
        );

    \I__9872\ : InMux
    port map (
            O => \N__43983\,
            I => \N__43974\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__43980\,
            I => \N__43969\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__43977\,
            I => \N__43969\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__43974\,
            I => \N__43965\
        );

    \I__9868\ : Span4Mux_v
    port map (
            O => \N__43969\,
            I => \N__43962\
        );

    \I__9867\ : InMux
    port map (
            O => \N__43968\,
            I => \N__43959\
        );

    \I__9866\ : Span4Mux_v
    port map (
            O => \N__43965\,
            I => \N__43956\
        );

    \I__9865\ : Span4Mux_h
    port map (
            O => \N__43962\,
            I => \N__43951\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__43959\,
            I => \N__43951\
        );

    \I__9863\ : Odrv4
    port map (
            O => \N__43956\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__9862\ : Odrv4
    port map (
            O => \N__43951\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__9861\ : InMux
    port map (
            O => \N__43946\,
            I => \bfn_18_10_0_\
        );

    \I__9860\ : CascadeMux
    port map (
            O => \N__43943\,
            I => \N__43939\
        );

    \I__9859\ : InMux
    port map (
            O => \N__43942\,
            I => \N__43936\
        );

    \I__9858\ : InMux
    port map (
            O => \N__43939\,
            I => \N__43932\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__43936\,
            I => \N__43929\
        );

    \I__9856\ : InMux
    port map (
            O => \N__43935\,
            I => \N__43926\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__43932\,
            I => \N__43923\
        );

    \I__9854\ : Span4Mux_h
    port map (
            O => \N__43929\,
            I => \N__43920\
        );

    \I__9853\ : LocalMux
    port map (
            O => \N__43926\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__9852\ : Odrv4
    port map (
            O => \N__43923\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__9851\ : Odrv4
    port map (
            O => \N__43920\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__9850\ : InMux
    port map (
            O => \N__43913\,
            I => \N__43906\
        );

    \I__9849\ : InMux
    port map (
            O => \N__43912\,
            I => \N__43906\
        );

    \I__9848\ : InMux
    port map (
            O => \N__43911\,
            I => \N__43902\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__43906\,
            I => \N__43899\
        );

    \I__9846\ : InMux
    port map (
            O => \N__43905\,
            I => \N__43896\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__43902\,
            I => \N__43893\
        );

    \I__9844\ : Span4Mux_h
    port map (
            O => \N__43899\,
            I => \N__43890\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__43896\,
            I => \N__43887\
        );

    \I__9842\ : Odrv4
    port map (
            O => \N__43893\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9841\ : Odrv4
    port map (
            O => \N__43890\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9840\ : Odrv4
    port map (
            O => \N__43887\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9839\ : InMux
    port map (
            O => \N__43880\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__9838\ : InMux
    port map (
            O => \N__43877\,
            I => \N__43870\
        );

    \I__9837\ : InMux
    port map (
            O => \N__43876\,
            I => \N__43870\
        );

    \I__9836\ : InMux
    port map (
            O => \N__43875\,
            I => \N__43867\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__43870\,
            I => \N__43864\
        );

    \I__9834\ : LocalMux
    port map (
            O => \N__43867\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__9833\ : Odrv4
    port map (
            O => \N__43864\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__9832\ : CascadeMux
    port map (
            O => \N__43859\,
            I => \N__43856\
        );

    \I__9831\ : InMux
    port map (
            O => \N__43856\,
            I => \N__43852\
        );

    \I__9830\ : InMux
    port map (
            O => \N__43855\,
            I => \N__43849\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__43852\,
            I => \N__43846\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__43849\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__9827\ : Odrv4
    port map (
            O => \N__43846\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__9826\ : InMux
    port map (
            O => \N__43841\,
            I => \N__43834\
        );

    \I__9825\ : InMux
    port map (
            O => \N__43840\,
            I => \N__43834\
        );

    \I__9824\ : InMux
    port map (
            O => \N__43839\,
            I => \N__43831\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__43834\,
            I => \N__43828\
        );

    \I__9822\ : LocalMux
    port map (
            O => \N__43831\,
            I => \N__43824\
        );

    \I__9821\ : Span4Mux_h
    port map (
            O => \N__43828\,
            I => \N__43821\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43827\,
            I => \N__43818\
        );

    \I__9819\ : Odrv4
    port map (
            O => \N__43824\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__9818\ : Odrv4
    port map (
            O => \N__43821\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__43818\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__9816\ : InMux
    port map (
            O => \N__43811\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__9815\ : InMux
    port map (
            O => \N__43808\,
            I => \N__43805\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__43805\,
            I => \N__43801\
        );

    \I__9813\ : InMux
    port map (
            O => \N__43804\,
            I => \N__43798\
        );

    \I__9812\ : Span4Mux_v
    port map (
            O => \N__43801\,
            I => \N__43795\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__43798\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__9810\ : Odrv4
    port map (
            O => \N__43795\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__9809\ : CascadeMux
    port map (
            O => \N__43790\,
            I => \N__43787\
        );

    \I__9808\ : InMux
    port map (
            O => \N__43787\,
            I => \N__43783\
        );

    \I__9807\ : InMux
    port map (
            O => \N__43786\,
            I => \N__43780\
        );

    \I__9806\ : LocalMux
    port map (
            O => \N__43783\,
            I => \N__43774\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__43780\,
            I => \N__43774\
        );

    \I__9804\ : InMux
    port map (
            O => \N__43779\,
            I => \N__43771\
        );

    \I__9803\ : Span4Mux_h
    port map (
            O => \N__43774\,
            I => \N__43768\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__43771\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__9801\ : Odrv4
    port map (
            O => \N__43768\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__9800\ : InMux
    port map (
            O => \N__43763\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__9799\ : InMux
    port map (
            O => \N__43760\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__9798\ : CascadeMux
    port map (
            O => \N__43757\,
            I => \N__43754\
        );

    \I__9797\ : InMux
    port map (
            O => \N__43754\,
            I => \N__43751\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__43751\,
            I => \N__43746\
        );

    \I__9795\ : InMux
    port map (
            O => \N__43750\,
            I => \N__43743\
        );

    \I__9794\ : InMux
    port map (
            O => \N__43749\,
            I => \N__43740\
        );

    \I__9793\ : Span4Mux_h
    port map (
            O => \N__43746\,
            I => \N__43737\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__43743\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9791\ : LocalMux
    port map (
            O => \N__43740\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9790\ : Odrv4
    port map (
            O => \N__43737\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9789\ : CascadeMux
    port map (
            O => \N__43730\,
            I => \N__43727\
        );

    \I__9788\ : InMux
    port map (
            O => \N__43727\,
            I => \N__43724\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__43724\,
            I => \N__43719\
        );

    \I__9786\ : InMux
    port map (
            O => \N__43723\,
            I => \N__43716\
        );

    \I__9785\ : InMux
    port map (
            O => \N__43722\,
            I => \N__43713\
        );

    \I__9784\ : Span12Mux_s8_h
    port map (
            O => \N__43719\,
            I => \N__43710\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__43716\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__43713\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__9781\ : Odrv12
    port map (
            O => \N__43710\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__9780\ : InMux
    port map (
            O => \N__43703\,
            I => \N__43697\
        );

    \I__9779\ : InMux
    port map (
            O => \N__43702\,
            I => \N__43694\
        );

    \I__9778\ : InMux
    port map (
            O => \N__43701\,
            I => \N__43691\
        );

    \I__9777\ : CascadeMux
    port map (
            O => \N__43700\,
            I => \N__43688\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__43697\,
            I => \N__43685\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__43694\,
            I => \N__43682\
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__43691\,
            I => \N__43679\
        );

    \I__9773\ : InMux
    port map (
            O => \N__43688\,
            I => \N__43676\
        );

    \I__9772\ : Span4Mux_h
    port map (
            O => \N__43685\,
            I => \N__43671\
        );

    \I__9771\ : Span4Mux_h
    port map (
            O => \N__43682\,
            I => \N__43671\
        );

    \I__9770\ : Span4Mux_h
    port map (
            O => \N__43679\,
            I => \N__43668\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__43676\,
            I => \N__43665\
        );

    \I__9768\ : Sp12to4
    port map (
            O => \N__43671\,
            I => \N__43662\
        );

    \I__9767\ : Span4Mux_v
    port map (
            O => \N__43668\,
            I => \N__43657\
        );

    \I__9766\ : Span4Mux_h
    port map (
            O => \N__43665\,
            I => \N__43657\
        );

    \I__9765\ : Odrv12
    port map (
            O => \N__43662\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__9764\ : Odrv4
    port map (
            O => \N__43657\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__9763\ : CEMux
    port map (
            O => \N__43652\,
            I => \N__43646\
        );

    \I__9762\ : CEMux
    port map (
            O => \N__43651\,
            I => \N__43642\
        );

    \I__9761\ : CEMux
    port map (
            O => \N__43650\,
            I => \N__43639\
        );

    \I__9760\ : CEMux
    port map (
            O => \N__43649\,
            I => \N__43636\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__43646\,
            I => \N__43633\
        );

    \I__9758\ : CEMux
    port map (
            O => \N__43645\,
            I => \N__43630\
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__43642\,
            I => \N__43627\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__43639\,
            I => \N__43624\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__43636\,
            I => \N__43621\
        );

    \I__9754\ : Span4Mux_h
    port map (
            O => \N__43633\,
            I => \N__43618\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__43630\,
            I => \N__43615\
        );

    \I__9752\ : Span4Mux_v
    port map (
            O => \N__43627\,
            I => \N__43612\
        );

    \I__9751\ : Span4Mux_v
    port map (
            O => \N__43624\,
            I => \N__43609\
        );

    \I__9750\ : Span4Mux_v
    port map (
            O => \N__43621\,
            I => \N__43606\
        );

    \I__9749\ : Span4Mux_h
    port map (
            O => \N__43618\,
            I => \N__43603\
        );

    \I__9748\ : Span4Mux_h
    port map (
            O => \N__43615\,
            I => \N__43600\
        );

    \I__9747\ : Span4Mux_h
    port map (
            O => \N__43612\,
            I => \N__43595\
        );

    \I__9746\ : Span4Mux_h
    port map (
            O => \N__43609\,
            I => \N__43595\
        );

    \I__9745\ : Span4Mux_h
    port map (
            O => \N__43606\,
            I => \N__43592\
        );

    \I__9744\ : Span4Mux_v
    port map (
            O => \N__43603\,
            I => \N__43587\
        );

    \I__9743\ : Span4Mux_h
    port map (
            O => \N__43600\,
            I => \N__43587\
        );

    \I__9742\ : Odrv4
    port map (
            O => \N__43595\,
            I => \delay_measurement_inst.delay_hc_timer.N_163_i\
        );

    \I__9741\ : Odrv4
    port map (
            O => \N__43592\,
            I => \delay_measurement_inst.delay_hc_timer.N_163_i\
        );

    \I__9740\ : Odrv4
    port map (
            O => \N__43587\,
            I => \delay_measurement_inst.delay_hc_timer.N_163_i\
        );

    \I__9739\ : InMux
    port map (
            O => \N__43580\,
            I => \N__43574\
        );

    \I__9738\ : InMux
    port map (
            O => \N__43579\,
            I => \N__43574\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__43574\,
            I => \N__43570\
        );

    \I__9736\ : InMux
    port map (
            O => \N__43573\,
            I => \N__43567\
        );

    \I__9735\ : Span4Mux_h
    port map (
            O => \N__43570\,
            I => \N__43564\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__43567\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__9733\ : Odrv4
    port map (
            O => \N__43564\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__9732\ : InMux
    port map (
            O => \N__43559\,
            I => \N__43556\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__43556\,
            I => \N__43551\
        );

    \I__9730\ : InMux
    port map (
            O => \N__43555\,
            I => \N__43548\
        );

    \I__9729\ : InMux
    port map (
            O => \N__43554\,
            I => \N__43545\
        );

    \I__9728\ : Span4Mux_h
    port map (
            O => \N__43551\,
            I => \N__43541\
        );

    \I__9727\ : LocalMux
    port map (
            O => \N__43548\,
            I => \N__43536\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__43545\,
            I => \N__43536\
        );

    \I__9725\ : InMux
    port map (
            O => \N__43544\,
            I => \N__43533\
        );

    \I__9724\ : Odrv4
    port map (
            O => \N__43541\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__9723\ : Odrv12
    port map (
            O => \N__43536\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__43533\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__9721\ : InMux
    port map (
            O => \N__43526\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__9720\ : CascadeMux
    port map (
            O => \N__43523\,
            I => \N__43520\
        );

    \I__9719\ : InMux
    port map (
            O => \N__43520\,
            I => \N__43516\
        );

    \I__9718\ : InMux
    port map (
            O => \N__43519\,
            I => \N__43513\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__43516\,
            I => \N__43509\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__43513\,
            I => \N__43506\
        );

    \I__9715\ : InMux
    port map (
            O => \N__43512\,
            I => \N__43503\
        );

    \I__9714\ : Span4Mux_h
    port map (
            O => \N__43509\,
            I => \N__43500\
        );

    \I__9713\ : Span4Mux_h
    port map (
            O => \N__43506\,
            I => \N__43497\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__43503\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__9711\ : Odrv4
    port map (
            O => \N__43500\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__9710\ : Odrv4
    port map (
            O => \N__43497\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__9709\ : InMux
    port map (
            O => \N__43490\,
            I => \N__43483\
        );

    \I__9708\ : InMux
    port map (
            O => \N__43489\,
            I => \N__43483\
        );

    \I__9707\ : InMux
    port map (
            O => \N__43488\,
            I => \N__43480\
        );

    \I__9706\ : LocalMux
    port map (
            O => \N__43483\,
            I => \N__43477\
        );

    \I__9705\ : LocalMux
    port map (
            O => \N__43480\,
            I => \N__43471\
        );

    \I__9704\ : Span12Mux_s8_v
    port map (
            O => \N__43477\,
            I => \N__43471\
        );

    \I__9703\ : InMux
    port map (
            O => \N__43476\,
            I => \N__43468\
        );

    \I__9702\ : Odrv12
    port map (
            O => \N__43471\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__9701\ : LocalMux
    port map (
            O => \N__43468\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__9700\ : InMux
    port map (
            O => \N__43463\,
            I => \bfn_18_9_0_\
        );

    \I__9699\ : CascadeMux
    port map (
            O => \N__43460\,
            I => \N__43456\
        );

    \I__9698\ : CascadeMux
    port map (
            O => \N__43459\,
            I => \N__43453\
        );

    \I__9697\ : InMux
    port map (
            O => \N__43456\,
            I => \N__43450\
        );

    \I__9696\ : InMux
    port map (
            O => \N__43453\,
            I => \N__43446\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__43450\,
            I => \N__43443\
        );

    \I__9694\ : InMux
    port map (
            O => \N__43449\,
            I => \N__43440\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__43446\,
            I => \N__43437\
        );

    \I__9692\ : Span4Mux_h
    port map (
            O => \N__43443\,
            I => \N__43434\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__43440\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__9690\ : Odrv4
    port map (
            O => \N__43437\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__9689\ : Odrv4
    port map (
            O => \N__43434\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__9688\ : InMux
    port map (
            O => \N__43427\,
            I => \N__43422\
        );

    \I__9687\ : InMux
    port map (
            O => \N__43426\,
            I => \N__43417\
        );

    \I__9686\ : InMux
    port map (
            O => \N__43425\,
            I => \N__43417\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__43422\,
            I => \N__43413\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__43417\,
            I => \N__43410\
        );

    \I__9683\ : CascadeMux
    port map (
            O => \N__43416\,
            I => \N__43407\
        );

    \I__9682\ : Span4Mux_h
    port map (
            O => \N__43413\,
            I => \N__43404\
        );

    \I__9681\ : Span12Mux_s8_v
    port map (
            O => \N__43410\,
            I => \N__43401\
        );

    \I__9680\ : InMux
    port map (
            O => \N__43407\,
            I => \N__43398\
        );

    \I__9679\ : Odrv4
    port map (
            O => \N__43404\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9678\ : Odrv12
    port map (
            O => \N__43401\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__43398\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9676\ : InMux
    port map (
            O => \N__43391\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__9675\ : InMux
    port map (
            O => \N__43388\,
            I => \N__43381\
        );

    \I__9674\ : InMux
    port map (
            O => \N__43387\,
            I => \N__43381\
        );

    \I__9673\ : InMux
    port map (
            O => \N__43386\,
            I => \N__43378\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__43381\,
            I => \N__43375\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__43378\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__9670\ : Odrv4
    port map (
            O => \N__43375\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__9669\ : InMux
    port map (
            O => \N__43370\,
            I => \N__43365\
        );

    \I__9668\ : InMux
    port map (
            O => \N__43369\,
            I => \N__43362\
        );

    \I__9667\ : InMux
    port map (
            O => \N__43368\,
            I => \N__43359\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__43365\,
            I => \N__43356\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__43362\,
            I => \N__43351\
        );

    \I__9664\ : LocalMux
    port map (
            O => \N__43359\,
            I => \N__43351\
        );

    \I__9663\ : Span4Mux_v
    port map (
            O => \N__43356\,
            I => \N__43347\
        );

    \I__9662\ : Span12Mux_s8_v
    port map (
            O => \N__43351\,
            I => \N__43344\
        );

    \I__9661\ : InMux
    port map (
            O => \N__43350\,
            I => \N__43341\
        );

    \I__9660\ : Odrv4
    port map (
            O => \N__43347\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__9659\ : Odrv12
    port map (
            O => \N__43344\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__43341\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__9657\ : InMux
    port map (
            O => \N__43334\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__9656\ : InMux
    port map (
            O => \N__43331\,
            I => \N__43324\
        );

    \I__9655\ : InMux
    port map (
            O => \N__43330\,
            I => \N__43324\
        );

    \I__9654\ : InMux
    port map (
            O => \N__43329\,
            I => \N__43321\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__43324\,
            I => \N__43318\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__43321\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__9651\ : Odrv4
    port map (
            O => \N__43318\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__9650\ : InMux
    port map (
            O => \N__43313\,
            I => \N__43310\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__43310\,
            I => \N__43305\
        );

    \I__9648\ : InMux
    port map (
            O => \N__43309\,
            I => \N__43300\
        );

    \I__9647\ : InMux
    port map (
            O => \N__43308\,
            I => \N__43300\
        );

    \I__9646\ : Span4Mux_v
    port map (
            O => \N__43305\,
            I => \N__43294\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__43300\,
            I => \N__43294\
        );

    \I__9644\ : CascadeMux
    port map (
            O => \N__43299\,
            I => \N__43291\
        );

    \I__9643\ : Span4Mux_v
    port map (
            O => \N__43294\,
            I => \N__43288\
        );

    \I__9642\ : InMux
    port map (
            O => \N__43291\,
            I => \N__43285\
        );

    \I__9641\ : Odrv4
    port map (
            O => \N__43288\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__43285\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9639\ : InMux
    port map (
            O => \N__43280\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__9638\ : CascadeMux
    port map (
            O => \N__43277\,
            I => \N__43273\
        );

    \I__9637\ : CascadeMux
    port map (
            O => \N__43276\,
            I => \N__43270\
        );

    \I__9636\ : InMux
    port map (
            O => \N__43273\,
            I => \N__43264\
        );

    \I__9635\ : InMux
    port map (
            O => \N__43270\,
            I => \N__43264\
        );

    \I__9634\ : InMux
    port map (
            O => \N__43269\,
            I => \N__43261\
        );

    \I__9633\ : LocalMux
    port map (
            O => \N__43264\,
            I => \N__43258\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__43261\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__9631\ : Odrv4
    port map (
            O => \N__43258\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__9630\ : InMux
    port map (
            O => \N__43253\,
            I => \N__43248\
        );

    \I__9629\ : InMux
    port map (
            O => \N__43252\,
            I => \N__43243\
        );

    \I__9628\ : InMux
    port map (
            O => \N__43251\,
            I => \N__43243\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__43248\,
            I => \N__43240\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__43243\,
            I => \N__43237\
        );

    \I__9625\ : Span4Mux_h
    port map (
            O => \N__43240\,
            I => \N__43233\
        );

    \I__9624\ : Span4Mux_h
    port map (
            O => \N__43237\,
            I => \N__43230\
        );

    \I__9623\ : InMux
    port map (
            O => \N__43236\,
            I => \N__43227\
        );

    \I__9622\ : Odrv4
    port map (
            O => \N__43233\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9621\ : Odrv4
    port map (
            O => \N__43230\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9620\ : LocalMux
    port map (
            O => \N__43227\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9619\ : InMux
    port map (
            O => \N__43220\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__9618\ : CascadeMux
    port map (
            O => \N__43217\,
            I => \N__43213\
        );

    \I__9617\ : CascadeMux
    port map (
            O => \N__43216\,
            I => \N__43210\
        );

    \I__9616\ : InMux
    port map (
            O => \N__43213\,
            I => \N__43205\
        );

    \I__9615\ : InMux
    port map (
            O => \N__43210\,
            I => \N__43205\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__43205\,
            I => \N__43201\
        );

    \I__9613\ : InMux
    port map (
            O => \N__43204\,
            I => \N__43198\
        );

    \I__9612\ : Span4Mux_v
    port map (
            O => \N__43201\,
            I => \N__43195\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__43198\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__9610\ : Odrv4
    port map (
            O => \N__43195\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__9609\ : InMux
    port map (
            O => \N__43190\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__9608\ : CascadeMux
    port map (
            O => \N__43187\,
            I => \N__43184\
        );

    \I__9607\ : InMux
    port map (
            O => \N__43184\,
            I => \N__43180\
        );

    \I__9606\ : InMux
    port map (
            O => \N__43183\,
            I => \N__43177\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__43180\,
            I => \N__43171\
        );

    \I__9604\ : LocalMux
    port map (
            O => \N__43177\,
            I => \N__43171\
        );

    \I__9603\ : InMux
    port map (
            O => \N__43176\,
            I => \N__43168\
        );

    \I__9602\ : Span4Mux_h
    port map (
            O => \N__43171\,
            I => \N__43165\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__43168\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__9600\ : Odrv4
    port map (
            O => \N__43165\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__9599\ : InMux
    port map (
            O => \N__43160\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__9598\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43154\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__43154\,
            I => \N__43151\
        );

    \I__9596\ : Span4Mux_h
    port map (
            O => \N__43151\,
            I => \N__43147\
        );

    \I__9595\ : CascadeMux
    port map (
            O => \N__43150\,
            I => \N__43142\
        );

    \I__9594\ : Span4Mux_v
    port map (
            O => \N__43147\,
            I => \N__43139\
        );

    \I__9593\ : InMux
    port map (
            O => \N__43146\,
            I => \N__43134\
        );

    \I__9592\ : InMux
    port map (
            O => \N__43145\,
            I => \N__43134\
        );

    \I__9591\ : InMux
    port map (
            O => \N__43142\,
            I => \N__43131\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__43139\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__43134\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__43131\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__9587\ : InMux
    port map (
            O => \N__43124\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__9586\ : CascadeMux
    port map (
            O => \N__43121\,
            I => \N__43117\
        );

    \I__9585\ : CascadeMux
    port map (
            O => \N__43120\,
            I => \N__43114\
        );

    \I__9584\ : InMux
    port map (
            O => \N__43117\,
            I => \N__43111\
        );

    \I__9583\ : InMux
    port map (
            O => \N__43114\,
            I => \N__43108\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__43111\,
            I => \N__43104\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__43108\,
            I => \N__43101\
        );

    \I__9580\ : InMux
    port map (
            O => \N__43107\,
            I => \N__43098\
        );

    \I__9579\ : Span4Mux_h
    port map (
            O => \N__43104\,
            I => \N__43095\
        );

    \I__9578\ : Span4Mux_h
    port map (
            O => \N__43101\,
            I => \N__43092\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__43098\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9576\ : Odrv4
    port map (
            O => \N__43095\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9575\ : Odrv4
    port map (
            O => \N__43092\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9574\ : InMux
    port map (
            O => \N__43085\,
            I => \N__43082\
        );

    \I__9573\ : LocalMux
    port map (
            O => \N__43082\,
            I => \N__43079\
        );

    \I__9572\ : Span4Mux_v
    port map (
            O => \N__43079\,
            I => \N__43073\
        );

    \I__9571\ : InMux
    port map (
            O => \N__43078\,
            I => \N__43070\
        );

    \I__9570\ : InMux
    port map (
            O => \N__43077\,
            I => \N__43065\
        );

    \I__9569\ : InMux
    port map (
            O => \N__43076\,
            I => \N__43065\
        );

    \I__9568\ : Odrv4
    port map (
            O => \N__43073\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__43070\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__43065\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__9565\ : InMux
    port map (
            O => \N__43058\,
            I => \bfn_18_8_0_\
        );

    \I__9564\ : CascadeMux
    port map (
            O => \N__43055\,
            I => \N__43051\
        );

    \I__9563\ : InMux
    port map (
            O => \N__43054\,
            I => \N__43048\
        );

    \I__9562\ : InMux
    port map (
            O => \N__43051\,
            I => \N__43044\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__43048\,
            I => \N__43041\
        );

    \I__9560\ : InMux
    port map (
            O => \N__43047\,
            I => \N__43038\
        );

    \I__9559\ : LocalMux
    port map (
            O => \N__43044\,
            I => \N__43033\
        );

    \I__9558\ : Span4Mux_h
    port map (
            O => \N__43041\,
            I => \N__43033\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__43038\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__9556\ : Odrv4
    port map (
            O => \N__43033\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__9555\ : InMux
    port map (
            O => \N__43028\,
            I => \N__43025\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__43025\,
            I => \N__43021\
        );

    \I__9553\ : InMux
    port map (
            O => \N__43024\,
            I => \N__43018\
        );

    \I__9552\ : Span4Mux_v
    port map (
            O => \N__43021\,
            I => \N__43013\
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__43018\,
            I => \N__43010\
        );

    \I__9550\ : InMux
    port map (
            O => \N__43017\,
            I => \N__43005\
        );

    \I__9549\ : InMux
    port map (
            O => \N__43016\,
            I => \N__43005\
        );

    \I__9548\ : Odrv4
    port map (
            O => \N__43013\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__9547\ : Odrv4
    port map (
            O => \N__43010\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__43005\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__9545\ : InMux
    port map (
            O => \N__42998\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__9544\ : InMux
    port map (
            O => \N__42995\,
            I => \N__42988\
        );

    \I__9543\ : InMux
    port map (
            O => \N__42994\,
            I => \N__42988\
        );

    \I__9542\ : InMux
    port map (
            O => \N__42993\,
            I => \N__42985\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__42988\,
            I => \N__42982\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__42985\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__9539\ : Odrv4
    port map (
            O => \N__42982\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__9538\ : InMux
    port map (
            O => \N__42977\,
            I => \N__42974\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__42974\,
            I => \N__42968\
        );

    \I__9536\ : InMux
    port map (
            O => \N__42973\,
            I => \N__42963\
        );

    \I__9535\ : InMux
    port map (
            O => \N__42972\,
            I => \N__42963\
        );

    \I__9534\ : InMux
    port map (
            O => \N__42971\,
            I => \N__42960\
        );

    \I__9533\ : Odrv4
    port map (
            O => \N__42968\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__42963\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__42960\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__9530\ : InMux
    port map (
            O => \N__42953\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__9529\ : InMux
    port map (
            O => \N__42950\,
            I => \N__42943\
        );

    \I__9528\ : InMux
    port map (
            O => \N__42949\,
            I => \N__42943\
        );

    \I__9527\ : InMux
    port map (
            O => \N__42948\,
            I => \N__42940\
        );

    \I__9526\ : LocalMux
    port map (
            O => \N__42943\,
            I => \N__42937\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__42940\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__9524\ : Odrv4
    port map (
            O => \N__42937\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__9523\ : InMux
    port map (
            O => \N__42932\,
            I => \N__42929\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__42929\,
            I => \N__42924\
        );

    \I__9521\ : InMux
    port map (
            O => \N__42928\,
            I => \N__42921\
        );

    \I__9520\ : InMux
    port map (
            O => \N__42927\,
            I => \N__42918\
        );

    \I__9519\ : Span4Mux_h
    port map (
            O => \N__42924\,
            I => \N__42914\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__42921\,
            I => \N__42909\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__42918\,
            I => \N__42909\
        );

    \I__9516\ : InMux
    port map (
            O => \N__42917\,
            I => \N__42906\
        );

    \I__9515\ : Odrv4
    port map (
            O => \N__42914\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__9514\ : Odrv4
    port map (
            O => \N__42909\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__42906\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__9512\ : InMux
    port map (
            O => \N__42899\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__9511\ : CascadeMux
    port map (
            O => \N__42896\,
            I => \N__42892\
        );

    \I__9510\ : CascadeMux
    port map (
            O => \N__42895\,
            I => \N__42889\
        );

    \I__9509\ : InMux
    port map (
            O => \N__42892\,
            I => \N__42883\
        );

    \I__9508\ : InMux
    port map (
            O => \N__42889\,
            I => \N__42883\
        );

    \I__9507\ : InMux
    port map (
            O => \N__42888\,
            I => \N__42880\
        );

    \I__9506\ : LocalMux
    port map (
            O => \N__42883\,
            I => \N__42877\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__42880\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__9504\ : Odrv4
    port map (
            O => \N__42877\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__9503\ : InMux
    port map (
            O => \N__42872\,
            I => \N__42869\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__42869\,
            I => \N__42864\
        );

    \I__9501\ : InMux
    port map (
            O => \N__42868\,
            I => \N__42859\
        );

    \I__9500\ : InMux
    port map (
            O => \N__42867\,
            I => \N__42859\
        );

    \I__9499\ : Span4Mux_v
    port map (
            O => \N__42864\,
            I => \N__42855\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42859\,
            I => \N__42852\
        );

    \I__9497\ : InMux
    port map (
            O => \N__42858\,
            I => \N__42849\
        );

    \I__9496\ : Odrv4
    port map (
            O => \N__42855\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__9495\ : Odrv12
    port map (
            O => \N__42852\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__42849\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__9493\ : InMux
    port map (
            O => \N__42842\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__9492\ : CascadeMux
    port map (
            O => \N__42839\,
            I => \N__42835\
        );

    \I__9491\ : CascadeMux
    port map (
            O => \N__42838\,
            I => \N__42832\
        );

    \I__9490\ : InMux
    port map (
            O => \N__42835\,
            I => \N__42827\
        );

    \I__9489\ : InMux
    port map (
            O => \N__42832\,
            I => \N__42827\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__42827\,
            I => \N__42823\
        );

    \I__9487\ : InMux
    port map (
            O => \N__42826\,
            I => \N__42820\
        );

    \I__9486\ : Span4Mux_v
    port map (
            O => \N__42823\,
            I => \N__42817\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__42820\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__9484\ : Odrv4
    port map (
            O => \N__42817\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__9483\ : InMux
    port map (
            O => \N__42812\,
            I => \N__42808\
        );

    \I__9482\ : InMux
    port map (
            O => \N__42811\,
            I => \N__42805\
        );

    \I__9481\ : LocalMux
    port map (
            O => \N__42808\,
            I => \N__42800\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__42805\,
            I => \N__42797\
        );

    \I__9479\ : InMux
    port map (
            O => \N__42804\,
            I => \N__42794\
        );

    \I__9478\ : CascadeMux
    port map (
            O => \N__42803\,
            I => \N__42791\
        );

    \I__9477\ : Span4Mux_v
    port map (
            O => \N__42800\,
            I => \N__42788\
        );

    \I__9476\ : Span4Mux_h
    port map (
            O => \N__42797\,
            I => \N__42783\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__42794\,
            I => \N__42783\
        );

    \I__9474\ : InMux
    port map (
            O => \N__42791\,
            I => \N__42780\
        );

    \I__9473\ : Odrv4
    port map (
            O => \N__42788\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__9472\ : Odrv4
    port map (
            O => \N__42783\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__42780\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__9470\ : InMux
    port map (
            O => \N__42773\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__9469\ : CascadeMux
    port map (
            O => \N__42770\,
            I => \N__42767\
        );

    \I__9468\ : InMux
    port map (
            O => \N__42767\,
            I => \N__42763\
        );

    \I__9467\ : InMux
    port map (
            O => \N__42766\,
            I => \N__42760\
        );

    \I__9466\ : LocalMux
    port map (
            O => \N__42763\,
            I => \N__42754\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__42760\,
            I => \N__42754\
        );

    \I__9464\ : InMux
    port map (
            O => \N__42759\,
            I => \N__42751\
        );

    \I__9463\ : Span4Mux_h
    port map (
            O => \N__42754\,
            I => \N__42748\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__42751\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__9461\ : Odrv4
    port map (
            O => \N__42748\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__9460\ : InMux
    port map (
            O => \N__42743\,
            I => \N__42738\
        );

    \I__9459\ : InMux
    port map (
            O => \N__42742\,
            I => \N__42733\
        );

    \I__9458\ : InMux
    port map (
            O => \N__42741\,
            I => \N__42733\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__42738\,
            I => \N__42730\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__42733\,
            I => \N__42727\
        );

    \I__9455\ : Span4Mux_h
    port map (
            O => \N__42730\,
            I => \N__42721\
        );

    \I__9454\ : Span4Mux_h
    port map (
            O => \N__42727\,
            I => \N__42721\
        );

    \I__9453\ : InMux
    port map (
            O => \N__42726\,
            I => \N__42718\
        );

    \I__9452\ : Odrv4
    port map (
            O => \N__42721\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__42718\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__9450\ : InMux
    port map (
            O => \N__42713\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__9449\ : InMux
    port map (
            O => \N__42710\,
            I => \N__42706\
        );

    \I__9448\ : InMux
    port map (
            O => \N__42709\,
            I => \N__42702\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__42706\,
            I => \N__42699\
        );

    \I__9446\ : InMux
    port map (
            O => \N__42705\,
            I => \N__42696\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__42702\,
            I => \N__42691\
        );

    \I__9444\ : Span4Mux_v
    port map (
            O => \N__42699\,
            I => \N__42691\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__42696\,
            I => \N__42688\
        );

    \I__9442\ : Odrv4
    port map (
            O => \N__42691\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__9441\ : Odrv4
    port map (
            O => \N__42688\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__9440\ : InMux
    port map (
            O => \N__42683\,
            I => \N__42680\
        );

    \I__9439\ : LocalMux
    port map (
            O => \N__42680\,
            I => \N__42677\
        );

    \I__9438\ : Span4Mux_h
    port map (
            O => \N__42677\,
            I => \N__42674\
        );

    \I__9437\ : Odrv4
    port map (
            O => \N__42674\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__9436\ : InMux
    port map (
            O => \N__42671\,
            I => \N__42667\
        );

    \I__9435\ : InMux
    port map (
            O => \N__42670\,
            I => \N__42663\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__42667\,
            I => \N__42660\
        );

    \I__9433\ : InMux
    port map (
            O => \N__42666\,
            I => \N__42657\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__42663\,
            I => \N__42654\
        );

    \I__9431\ : Span4Mux_h
    port map (
            O => \N__42660\,
            I => \N__42649\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__42657\,
            I => \N__42649\
        );

    \I__9429\ : Span4Mux_h
    port map (
            O => \N__42654\,
            I => \N__42643\
        );

    \I__9428\ : Span4Mux_h
    port map (
            O => \N__42649\,
            I => \N__42643\
        );

    \I__9427\ : InMux
    port map (
            O => \N__42648\,
            I => \N__42640\
        );

    \I__9426\ : Odrv4
    port map (
            O => \N__42643\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__9425\ : LocalMux
    port map (
            O => \N__42640\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__9424\ : InMux
    port map (
            O => \N__42635\,
            I => \N__42632\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__42632\,
            I => \N__42627\
        );

    \I__9422\ : InMux
    port map (
            O => \N__42631\,
            I => \N__42624\
        );

    \I__9421\ : InMux
    port map (
            O => \N__42630\,
            I => \N__42621\
        );

    \I__9420\ : Span4Mux_v
    port map (
            O => \N__42627\,
            I => \N__42618\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__42624\,
            I => \N__42613\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__42621\,
            I => \N__42613\
        );

    \I__9417\ : Span4Mux_h
    port map (
            O => \N__42618\,
            I => \N__42607\
        );

    \I__9416\ : Span4Mux_h
    port map (
            O => \N__42613\,
            I => \N__42607\
        );

    \I__9415\ : InMux
    port map (
            O => \N__42612\,
            I => \N__42604\
        );

    \I__9414\ : Odrv4
    port map (
            O => \N__42607\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__42604\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__9412\ : InMux
    port map (
            O => \N__42599\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__9411\ : InMux
    port map (
            O => \N__42596\,
            I => \N__42589\
        );

    \I__9410\ : InMux
    port map (
            O => \N__42595\,
            I => \N__42589\
        );

    \I__9409\ : InMux
    port map (
            O => \N__42594\,
            I => \N__42586\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__42589\,
            I => \N__42583\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__42586\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9406\ : Odrv4
    port map (
            O => \N__42583\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9405\ : InMux
    port map (
            O => \N__42578\,
            I => \N__42575\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__42575\,
            I => \N__42570\
        );

    \I__9403\ : InMux
    port map (
            O => \N__42574\,
            I => \N__42565\
        );

    \I__9402\ : InMux
    port map (
            O => \N__42573\,
            I => \N__42565\
        );

    \I__9401\ : Span4Mux_v
    port map (
            O => \N__42570\,
            I => \N__42560\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__42565\,
            I => \N__42560\
        );

    \I__9399\ : Span4Mux_h
    port map (
            O => \N__42560\,
            I => \N__42557\
        );

    \I__9398\ : Span4Mux_h
    port map (
            O => \N__42557\,
            I => \N__42553\
        );

    \I__9397\ : InMux
    port map (
            O => \N__42556\,
            I => \N__42550\
        );

    \I__9396\ : Odrv4
    port map (
            O => \N__42553\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__42550\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__9394\ : InMux
    port map (
            O => \N__42545\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__9393\ : InMux
    port map (
            O => \N__42542\,
            I => \N__42535\
        );

    \I__9392\ : InMux
    port map (
            O => \N__42541\,
            I => \N__42535\
        );

    \I__9391\ : InMux
    port map (
            O => \N__42540\,
            I => \N__42532\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__42535\,
            I => \N__42529\
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__42532\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9388\ : Odrv4
    port map (
            O => \N__42529\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9387\ : InMux
    port map (
            O => \N__42524\,
            I => \N__42521\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__42521\,
            I => \N__42517\
        );

    \I__9385\ : InMux
    port map (
            O => \N__42520\,
            I => \N__42514\
        );

    \I__9384\ : Span4Mux_v
    port map (
            O => \N__42517\,
            I => \N__42510\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__42514\,
            I => \N__42507\
        );

    \I__9382\ : InMux
    port map (
            O => \N__42513\,
            I => \N__42504\
        );

    \I__9381\ : Span4Mux_h
    port map (
            O => \N__42510\,
            I => \N__42500\
        );

    \I__9380\ : Span4Mux_v
    port map (
            O => \N__42507\,
            I => \N__42497\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__42504\,
            I => \N__42494\
        );

    \I__9378\ : InMux
    port map (
            O => \N__42503\,
            I => \N__42491\
        );

    \I__9377\ : Odrv4
    port map (
            O => \N__42500\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__9376\ : Odrv4
    port map (
            O => \N__42497\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__9375\ : Odrv12
    port map (
            O => \N__42494\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__42491\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__9373\ : InMux
    port map (
            O => \N__42482\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__9372\ : CascadeMux
    port map (
            O => \N__42479\,
            I => \N__42475\
        );

    \I__9371\ : CascadeMux
    port map (
            O => \N__42478\,
            I => \N__42472\
        );

    \I__9370\ : InMux
    port map (
            O => \N__42475\,
            I => \N__42466\
        );

    \I__9369\ : InMux
    port map (
            O => \N__42472\,
            I => \N__42466\
        );

    \I__9368\ : InMux
    port map (
            O => \N__42471\,
            I => \N__42463\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__42466\,
            I => \N__42460\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__42463\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9365\ : Odrv4
    port map (
            O => \N__42460\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9364\ : InMux
    port map (
            O => \N__42455\,
            I => \N__42451\
        );

    \I__9363\ : InMux
    port map (
            O => \N__42454\,
            I => \N__42447\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__42451\,
            I => \N__42444\
        );

    \I__9361\ : InMux
    port map (
            O => \N__42450\,
            I => \N__42441\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__42447\,
            I => \N__42438\
        );

    \I__9359\ : Span4Mux_v
    port map (
            O => \N__42444\,
            I => \N__42433\
        );

    \I__9358\ : LocalMux
    port map (
            O => \N__42441\,
            I => \N__42433\
        );

    \I__9357\ : Span4Mux_v
    port map (
            O => \N__42438\,
            I => \N__42429\
        );

    \I__9356\ : Span4Mux_h
    port map (
            O => \N__42433\,
            I => \N__42426\
        );

    \I__9355\ : InMux
    port map (
            O => \N__42432\,
            I => \N__42423\
        );

    \I__9354\ : Odrv4
    port map (
            O => \N__42429\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__9353\ : Odrv4
    port map (
            O => \N__42426\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__42423\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__9351\ : InMux
    port map (
            O => \N__42416\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__9350\ : CascadeMux
    port map (
            O => \N__42413\,
            I => \N__42409\
        );

    \I__9349\ : CascadeMux
    port map (
            O => \N__42412\,
            I => \N__42406\
        );

    \I__9348\ : InMux
    port map (
            O => \N__42409\,
            I => \N__42400\
        );

    \I__9347\ : InMux
    port map (
            O => \N__42406\,
            I => \N__42400\
        );

    \I__9346\ : InMux
    port map (
            O => \N__42405\,
            I => \N__42397\
        );

    \I__9345\ : LocalMux
    port map (
            O => \N__42400\,
            I => \N__42394\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__42397\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9343\ : Odrv4
    port map (
            O => \N__42394\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9342\ : InMux
    port map (
            O => \N__42389\,
            I => \N__42385\
        );

    \I__9341\ : InMux
    port map (
            O => \N__42388\,
            I => \N__42381\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__42385\,
            I => \N__42378\
        );

    \I__9339\ : InMux
    port map (
            O => \N__42384\,
            I => \N__42375\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__42381\,
            I => \N__42372\
        );

    \I__9337\ : Span4Mux_h
    port map (
            O => \N__42378\,
            I => \N__42369\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__42375\,
            I => \N__42364\
        );

    \I__9335\ : Span4Mux_h
    port map (
            O => \N__42372\,
            I => \N__42364\
        );

    \I__9334\ : Span4Mux_h
    port map (
            O => \N__42369\,
            I => \N__42358\
        );

    \I__9333\ : Span4Mux_h
    port map (
            O => \N__42364\,
            I => \N__42358\
        );

    \I__9332\ : InMux
    port map (
            O => \N__42363\,
            I => \N__42355\
        );

    \I__9331\ : Odrv4
    port map (
            O => \N__42358\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__42355\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__9329\ : InMux
    port map (
            O => \N__42350\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__9328\ : InMux
    port map (
            O => \N__42347\,
            I => \N__42341\
        );

    \I__9327\ : InMux
    port map (
            O => \N__42346\,
            I => \N__42341\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__42341\,
            I => \N__42337\
        );

    \I__9325\ : InMux
    port map (
            O => \N__42340\,
            I => \N__42334\
        );

    \I__9324\ : Span4Mux_h
    port map (
            O => \N__42337\,
            I => \N__42331\
        );

    \I__9323\ : LocalMux
    port map (
            O => \N__42334\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9322\ : Odrv4
    port map (
            O => \N__42331\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9321\ : InMux
    port map (
            O => \N__42326\,
            I => \N__42323\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__42323\,
            I => \N__42319\
        );

    \I__9319\ : InMux
    port map (
            O => \N__42322\,
            I => \N__42314\
        );

    \I__9318\ : Span4Mux_v
    port map (
            O => \N__42319\,
            I => \N__42311\
        );

    \I__9317\ : InMux
    port map (
            O => \N__42318\,
            I => \N__42308\
        );

    \I__9316\ : InMux
    port map (
            O => \N__42317\,
            I => \N__42305\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__42314\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__9314\ : Odrv4
    port map (
            O => \N__42311\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__42308\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__42305\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__9311\ : InMux
    port map (
            O => \N__42296\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__9310\ : CascadeMux
    port map (
            O => \N__42293\,
            I => \N__42290\
        );

    \I__9309\ : InMux
    port map (
            O => \N__42290\,
            I => \N__42286\
        );

    \I__9308\ : InMux
    port map (
            O => \N__42289\,
            I => \N__42283\
        );

    \I__9307\ : LocalMux
    port map (
            O => \N__42286\,
            I => \N__42277\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__42283\,
            I => \N__42277\
        );

    \I__9305\ : InMux
    port map (
            O => \N__42282\,
            I => \N__42274\
        );

    \I__9304\ : Span4Mux_h
    port map (
            O => \N__42277\,
            I => \N__42271\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__42274\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__9302\ : Odrv4
    port map (
            O => \N__42271\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__9301\ : InMux
    port map (
            O => \N__42266\,
            I => \N__42263\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__42263\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__9299\ : InMux
    port map (
            O => \N__42260\,
            I => \N__42257\
        );

    \I__9298\ : LocalMux
    port map (
            O => \N__42257\,
            I => \N__42254\
        );

    \I__9297\ : Odrv4
    port map (
            O => \N__42254\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__9296\ : InMux
    port map (
            O => \N__42251\,
            I => \N__42248\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__42248\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__9294\ : InMux
    port map (
            O => \N__42245\,
            I => \N__42242\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__42242\,
            I => \N__42239\
        );

    \I__9292\ : Odrv4
    port map (
            O => \N__42239\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__9291\ : InMux
    port map (
            O => \N__42236\,
            I => \N__42233\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__42233\,
            I => \N__42230\
        );

    \I__9289\ : Odrv4
    port map (
            O => \N__42230\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__9288\ : InMux
    port map (
            O => \N__42227\,
            I => \N__42224\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__42224\,
            I => \N__42221\
        );

    \I__9286\ : Span4Mux_v
    port map (
            O => \N__42221\,
            I => \N__42218\
        );

    \I__9285\ : Odrv4
    port map (
            O => \N__42218\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__9284\ : InMux
    port map (
            O => \N__42215\,
            I => \N__42212\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__42212\,
            I => \N__42209\
        );

    \I__9282\ : Odrv4
    port map (
            O => \N__42209\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__9281\ : InMux
    port map (
            O => \N__42206\,
            I => \N__42203\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__42203\,
            I => \N__42200\
        );

    \I__9279\ : Odrv4
    port map (
            O => \N__42200\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__9278\ : CascadeMux
    port map (
            O => \N__42197\,
            I => \N__42194\
        );

    \I__9277\ : InMux
    port map (
            O => \N__42194\,
            I => \N__42191\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__42191\,
            I => \N__42188\
        );

    \I__9275\ : Odrv4
    port map (
            O => \N__42188\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__9274\ : CascadeMux
    port map (
            O => \N__42185\,
            I => \N__42182\
        );

    \I__9273\ : InMux
    port map (
            O => \N__42182\,
            I => \N__42179\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__42179\,
            I => \N__42174\
        );

    \I__9271\ : InMux
    port map (
            O => \N__42178\,
            I => \N__42171\
        );

    \I__9270\ : InMux
    port map (
            O => \N__42177\,
            I => \N__42168\
        );

    \I__9269\ : Odrv12
    port map (
            O => \N__42174\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__42171\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__42168\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9266\ : CascadeMux
    port map (
            O => \N__42161\,
            I => \N__42158\
        );

    \I__9265\ : InMux
    port map (
            O => \N__42158\,
            I => \N__42155\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__42155\,
            I => \N__42152\
        );

    \I__9263\ : Odrv4
    port map (
            O => \N__42152\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__9262\ : CascadeMux
    port map (
            O => \N__42149\,
            I => \N__42146\
        );

    \I__9261\ : InMux
    port map (
            O => \N__42146\,
            I => \N__42143\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__42143\,
            I => \N__42140\
        );

    \I__9259\ : Odrv4
    port map (
            O => \N__42140\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__9258\ : InMux
    port map (
            O => \N__42137\,
            I => \N__42134\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__42134\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__9256\ : CascadeMux
    port map (
            O => \N__42131\,
            I => \N__42128\
        );

    \I__9255\ : InMux
    port map (
            O => \N__42128\,
            I => \N__42125\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__42125\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__9253\ : InMux
    port map (
            O => \N__42122\,
            I => \N__42119\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__42119\,
            I => \N__42116\
        );

    \I__9251\ : Odrv12
    port map (
            O => \N__42116\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__9250\ : InMux
    port map (
            O => \N__42113\,
            I => \N__42110\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__42110\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__9248\ : InMux
    port map (
            O => \N__42107\,
            I => \N__42104\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__42104\,
            I => \N__42101\
        );

    \I__9246\ : Odrv4
    port map (
            O => \N__42101\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__9245\ : InMux
    port map (
            O => \N__42098\,
            I => \N__42095\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__42095\,
            I => \N__42092\
        );

    \I__9243\ : Odrv4
    port map (
            O => \N__42092\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__9242\ : InMux
    port map (
            O => \N__42089\,
            I => \N__42086\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__42086\,
            I => \N__42083\
        );

    \I__9240\ : Odrv4
    port map (
            O => \N__42083\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__9239\ : InMux
    port map (
            O => \N__42080\,
            I => \N__42075\
        );

    \I__9238\ : InMux
    port map (
            O => \N__42079\,
            I => \N__42072\
        );

    \I__9237\ : InMux
    port map (
            O => \N__42078\,
            I => \N__42069\
        );

    \I__9236\ : LocalMux
    port map (
            O => \N__42075\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__42072\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__42069\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9233\ : InMux
    port map (
            O => \N__42062\,
            I => \N__42059\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__42059\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__9231\ : InMux
    port map (
            O => \N__42056\,
            I => \N__42053\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__42053\,
            I => \N__42048\
        );

    \I__9229\ : InMux
    port map (
            O => \N__42052\,
            I => \N__42045\
        );

    \I__9228\ : InMux
    port map (
            O => \N__42051\,
            I => \N__42042\
        );

    \I__9227\ : Odrv4
    port map (
            O => \N__42048\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__42045\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9225\ : LocalMux
    port map (
            O => \N__42042\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9224\ : CascadeMux
    port map (
            O => \N__42035\,
            I => \N__42032\
        );

    \I__9223\ : InMux
    port map (
            O => \N__42032\,
            I => \N__42029\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__42029\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__9221\ : InMux
    port map (
            O => \N__42026\,
            I => \N__42023\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__42023\,
            I => \N__42018\
        );

    \I__9219\ : CascadeMux
    port map (
            O => \N__42022\,
            I => \N__42015\
        );

    \I__9218\ : InMux
    port map (
            O => \N__42021\,
            I => \N__42012\
        );

    \I__9217\ : Span4Mux_v
    port map (
            O => \N__42018\,
            I => \N__42009\
        );

    \I__9216\ : InMux
    port map (
            O => \N__42015\,
            I => \N__42006\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__42012\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9214\ : Odrv4
    port map (
            O => \N__42009\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__42006\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9212\ : CascadeMux
    port map (
            O => \N__41999\,
            I => \N__41996\
        );

    \I__9211\ : InMux
    port map (
            O => \N__41996\,
            I => \N__41993\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__41993\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__9209\ : InMux
    port map (
            O => \N__41990\,
            I => \N__41987\
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__41987\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__9207\ : CascadeMux
    port map (
            O => \N__41984\,
            I => \N__41979\
        );

    \I__9206\ : InMux
    port map (
            O => \N__41983\,
            I => \N__41976\
        );

    \I__9205\ : InMux
    port map (
            O => \N__41982\,
            I => \N__41973\
        );

    \I__9204\ : InMux
    port map (
            O => \N__41979\,
            I => \N__41970\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__41976\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__41973\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__41970\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9200\ : InMux
    port map (
            O => \N__41963\,
            I => \N__41960\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__41960\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__9198\ : InMux
    port map (
            O => \N__41957\,
            I => \N__41954\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__41954\,
            I => \N__41951\
        );

    \I__9196\ : Odrv4
    port map (
            O => \N__41951\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__9195\ : InMux
    port map (
            O => \N__41948\,
            I => \N__41943\
        );

    \I__9194\ : InMux
    port map (
            O => \N__41947\,
            I => \N__41940\
        );

    \I__9193\ : InMux
    port map (
            O => \N__41946\,
            I => \N__41937\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__41943\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__41940\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__41937\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9189\ : InMux
    port map (
            O => \N__41930\,
            I => \N__41927\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__41927\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__9187\ : CascadeMux
    port map (
            O => \N__41924\,
            I => \N__41921\
        );

    \I__9186\ : InMux
    port map (
            O => \N__41921\,
            I => \N__41918\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__41918\,
            I => \N__41913\
        );

    \I__9184\ : InMux
    port map (
            O => \N__41917\,
            I => \N__41910\
        );

    \I__9183\ : InMux
    port map (
            O => \N__41916\,
            I => \N__41907\
        );

    \I__9182\ : Odrv4
    port map (
            O => \N__41913\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__41910\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__41907\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9179\ : CascadeMux
    port map (
            O => \N__41900\,
            I => \N__41897\
        );

    \I__9178\ : InMux
    port map (
            O => \N__41897\,
            I => \N__41894\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__41894\,
            I => \N__41891\
        );

    \I__9176\ : Odrv4
    port map (
            O => \N__41891\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__9175\ : CascadeMux
    port map (
            O => \N__41888\,
            I => \N__41885\
        );

    \I__9174\ : InMux
    port map (
            O => \N__41885\,
            I => \N__41882\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__41882\,
            I => \N__41879\
        );

    \I__9172\ : Odrv4
    port map (
            O => \N__41879\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__9171\ : InMux
    port map (
            O => \N__41876\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__9170\ : InMux
    port map (
            O => \N__41873\,
            I => \N__41858\
        );

    \I__9169\ : InMux
    port map (
            O => \N__41872\,
            I => \N__41855\
        );

    \I__9168\ : InMux
    port map (
            O => \N__41871\,
            I => \N__41838\
        );

    \I__9167\ : InMux
    port map (
            O => \N__41870\,
            I => \N__41838\
        );

    \I__9166\ : InMux
    port map (
            O => \N__41869\,
            I => \N__41838\
        );

    \I__9165\ : InMux
    port map (
            O => \N__41868\,
            I => \N__41838\
        );

    \I__9164\ : InMux
    port map (
            O => \N__41867\,
            I => \N__41838\
        );

    \I__9163\ : InMux
    port map (
            O => \N__41866\,
            I => \N__41838\
        );

    \I__9162\ : InMux
    port map (
            O => \N__41865\,
            I => \N__41838\
        );

    \I__9161\ : InMux
    port map (
            O => \N__41864\,
            I => \N__41838\
        );

    \I__9160\ : CascadeMux
    port map (
            O => \N__41863\,
            I => \N__41834\
        );

    \I__9159\ : InMux
    port map (
            O => \N__41862\,
            I => \N__41831\
        );

    \I__9158\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41828\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__41858\,
            I => \N__41815\
        );

    \I__9156\ : LocalMux
    port map (
            O => \N__41855\,
            I => \N__41815\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__41838\,
            I => \N__41815\
        );

    \I__9154\ : InMux
    port map (
            O => \N__41837\,
            I => \N__41812\
        );

    \I__9153\ : InMux
    port map (
            O => \N__41834\,
            I => \N__41797\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__41831\,
            I => \N__41792\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__41828\,
            I => \N__41792\
        );

    \I__9150\ : InMux
    port map (
            O => \N__41827\,
            I => \N__41789\
        );

    \I__9149\ : InMux
    port map (
            O => \N__41826\,
            I => \N__41778\
        );

    \I__9148\ : InMux
    port map (
            O => \N__41825\,
            I => \N__41778\
        );

    \I__9147\ : InMux
    port map (
            O => \N__41824\,
            I => \N__41778\
        );

    \I__9146\ : InMux
    port map (
            O => \N__41823\,
            I => \N__41778\
        );

    \I__9145\ : InMux
    port map (
            O => \N__41822\,
            I => \N__41778\
        );

    \I__9144\ : Span4Mux_v
    port map (
            O => \N__41815\,
            I => \N__41773\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__41812\,
            I => \N__41773\
        );

    \I__9142\ : InMux
    port map (
            O => \N__41811\,
            I => \N__41756\
        );

    \I__9141\ : InMux
    port map (
            O => \N__41810\,
            I => \N__41756\
        );

    \I__9140\ : InMux
    port map (
            O => \N__41809\,
            I => \N__41756\
        );

    \I__9139\ : InMux
    port map (
            O => \N__41808\,
            I => \N__41756\
        );

    \I__9138\ : InMux
    port map (
            O => \N__41807\,
            I => \N__41756\
        );

    \I__9137\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41756\
        );

    \I__9136\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41756\
        );

    \I__9135\ : InMux
    port map (
            O => \N__41804\,
            I => \N__41756\
        );

    \I__9134\ : InMux
    port map (
            O => \N__41803\,
            I => \N__41747\
        );

    \I__9133\ : InMux
    port map (
            O => \N__41802\,
            I => \N__41747\
        );

    \I__9132\ : InMux
    port map (
            O => \N__41801\,
            I => \N__41747\
        );

    \I__9131\ : InMux
    port map (
            O => \N__41800\,
            I => \N__41747\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__41797\,
            I => \N__41744\
        );

    \I__9129\ : Span4Mux_v
    port map (
            O => \N__41792\,
            I => \N__41737\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__41789\,
            I => \N__41737\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__41778\,
            I => \N__41737\
        );

    \I__9126\ : Span4Mux_h
    port map (
            O => \N__41773\,
            I => \N__41734\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__41756\,
            I => \N__41729\
        );

    \I__9124\ : LocalMux
    port map (
            O => \N__41747\,
            I => \N__41729\
        );

    \I__9123\ : Odrv4
    port map (
            O => \N__41744\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__9122\ : Odrv4
    port map (
            O => \N__41737\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__9121\ : Odrv4
    port map (
            O => \N__41734\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__9120\ : Odrv12
    port map (
            O => \N__41729\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__9119\ : InMux
    port map (
            O => \N__41720\,
            I => \N__41717\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__41717\,
            I => \N__41712\
        );

    \I__9117\ : InMux
    port map (
            O => \N__41716\,
            I => \N__41709\
        );

    \I__9116\ : InMux
    port map (
            O => \N__41715\,
            I => \N__41706\
        );

    \I__9115\ : Odrv4
    port map (
            O => \N__41712\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__41709\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__41706\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9112\ : CascadeMux
    port map (
            O => \N__41699\,
            I => \N__41696\
        );

    \I__9111\ : InMux
    port map (
            O => \N__41696\,
            I => \N__41693\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__41693\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__9109\ : InMux
    port map (
            O => \N__41690\,
            I => \N__41687\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__41687\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__9107\ : InMux
    port map (
            O => \N__41684\,
            I => \N__41681\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__41681\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__9105\ : CascadeMux
    port map (
            O => \N__41678\,
            I => \N__41675\
        );

    \I__9104\ : InMux
    port map (
            O => \N__41675\,
            I => \N__41672\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__41672\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__9102\ : CascadeMux
    port map (
            O => \N__41669\,
            I => \N__41666\
        );

    \I__9101\ : InMux
    port map (
            O => \N__41666\,
            I => \N__41663\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__41663\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__9099\ : CascadeMux
    port map (
            O => \N__41660\,
            I => \N__41657\
        );

    \I__9098\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41654\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__41654\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__9096\ : CascadeMux
    port map (
            O => \N__41651\,
            I => \N__41648\
        );

    \I__9095\ : InMux
    port map (
            O => \N__41648\,
            I => \N__41645\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41645\,
            I => \N__41642\
        );

    \I__9093\ : Span4Mux_h
    port map (
            O => \N__41642\,
            I => \N__41639\
        );

    \I__9092\ : Odrv4
    port map (
            O => \N__41639\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\
        );

    \I__9091\ : CascadeMux
    port map (
            O => \N__41636\,
            I => \N__41633\
        );

    \I__9090\ : InMux
    port map (
            O => \N__41633\,
            I => \N__41630\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__41630\,
            I => \N__41627\
        );

    \I__9088\ : Odrv4
    port map (
            O => \N__41627\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\
        );

    \I__9087\ : InMux
    port map (
            O => \N__41624\,
            I => \N__41621\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__41621\,
            I => \N__41618\
        );

    \I__9085\ : Span4Mux_h
    port map (
            O => \N__41618\,
            I => \N__41615\
        );

    \I__9084\ : Odrv4
    port map (
            O => \N__41615\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__9083\ : CascadeMux
    port map (
            O => \N__41612\,
            I => \N__41609\
        );

    \I__9082\ : InMux
    port map (
            O => \N__41609\,
            I => \N__41606\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__41606\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__9080\ : InMux
    port map (
            O => \N__41603\,
            I => \N__41600\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__41600\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__9078\ : CascadeMux
    port map (
            O => \N__41597\,
            I => \N__41594\
        );

    \I__9077\ : InMux
    port map (
            O => \N__41594\,
            I => \N__41591\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__41591\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__9075\ : InMux
    port map (
            O => \N__41588\,
            I => \N__41585\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__41585\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__9073\ : CascadeMux
    port map (
            O => \N__41582\,
            I => \N__41579\
        );

    \I__9072\ : InMux
    port map (
            O => \N__41579\,
            I => \N__41576\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__41576\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__9070\ : InMux
    port map (
            O => \N__41573\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__9069\ : InMux
    port map (
            O => \N__41570\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__9068\ : InMux
    port map (
            O => \N__41567\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__9067\ : InMux
    port map (
            O => \N__41564\,
            I => \N__41526\
        );

    \I__9066\ : InMux
    port map (
            O => \N__41563\,
            I => \N__41526\
        );

    \I__9065\ : InMux
    port map (
            O => \N__41562\,
            I => \N__41526\
        );

    \I__9064\ : InMux
    port map (
            O => \N__41561\,
            I => \N__41526\
        );

    \I__9063\ : InMux
    port map (
            O => \N__41560\,
            I => \N__41517\
        );

    \I__9062\ : InMux
    port map (
            O => \N__41559\,
            I => \N__41517\
        );

    \I__9061\ : InMux
    port map (
            O => \N__41558\,
            I => \N__41517\
        );

    \I__9060\ : InMux
    port map (
            O => \N__41557\,
            I => \N__41517\
        );

    \I__9059\ : InMux
    port map (
            O => \N__41556\,
            I => \N__41508\
        );

    \I__9058\ : InMux
    port map (
            O => \N__41555\,
            I => \N__41508\
        );

    \I__9057\ : InMux
    port map (
            O => \N__41554\,
            I => \N__41508\
        );

    \I__9056\ : InMux
    port map (
            O => \N__41553\,
            I => \N__41508\
        );

    \I__9055\ : InMux
    port map (
            O => \N__41552\,
            I => \N__41499\
        );

    \I__9054\ : InMux
    port map (
            O => \N__41551\,
            I => \N__41499\
        );

    \I__9053\ : InMux
    port map (
            O => \N__41550\,
            I => \N__41499\
        );

    \I__9052\ : InMux
    port map (
            O => \N__41549\,
            I => \N__41499\
        );

    \I__9051\ : InMux
    port map (
            O => \N__41548\,
            I => \N__41490\
        );

    \I__9050\ : InMux
    port map (
            O => \N__41547\,
            I => \N__41490\
        );

    \I__9049\ : InMux
    port map (
            O => \N__41546\,
            I => \N__41490\
        );

    \I__9048\ : InMux
    port map (
            O => \N__41545\,
            I => \N__41490\
        );

    \I__9047\ : InMux
    port map (
            O => \N__41544\,
            I => \N__41481\
        );

    \I__9046\ : InMux
    port map (
            O => \N__41543\,
            I => \N__41481\
        );

    \I__9045\ : InMux
    port map (
            O => \N__41542\,
            I => \N__41481\
        );

    \I__9044\ : InMux
    port map (
            O => \N__41541\,
            I => \N__41481\
        );

    \I__9043\ : InMux
    port map (
            O => \N__41540\,
            I => \N__41476\
        );

    \I__9042\ : InMux
    port map (
            O => \N__41539\,
            I => \N__41476\
        );

    \I__9041\ : InMux
    port map (
            O => \N__41538\,
            I => \N__41467\
        );

    \I__9040\ : InMux
    port map (
            O => \N__41537\,
            I => \N__41467\
        );

    \I__9039\ : InMux
    port map (
            O => \N__41536\,
            I => \N__41467\
        );

    \I__9038\ : InMux
    port map (
            O => \N__41535\,
            I => \N__41467\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__41526\,
            I => \N__41462\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__41517\,
            I => \N__41462\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__41508\,
            I => \N__41459\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__41499\,
            I => \N__41448\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__41490\,
            I => \N__41448\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__41481\,
            I => \N__41448\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__41476\,
            I => \N__41448\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__41467\,
            I => \N__41448\
        );

    \I__9029\ : Span4Mux_v
    port map (
            O => \N__41462\,
            I => \N__41441\
        );

    \I__9028\ : Span4Mux_h
    port map (
            O => \N__41459\,
            I => \N__41441\
        );

    \I__9027\ : Span4Mux_v
    port map (
            O => \N__41448\,
            I => \N__41441\
        );

    \I__9026\ : Span4Mux_h
    port map (
            O => \N__41441\,
            I => \N__41438\
        );

    \I__9025\ : Odrv4
    port map (
            O => \N__41438\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__9024\ : InMux
    port map (
            O => \N__41435\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__9023\ : CEMux
    port map (
            O => \N__41432\,
            I => \N__41427\
        );

    \I__9022\ : CEMux
    port map (
            O => \N__41431\,
            I => \N__41424\
        );

    \I__9021\ : CEMux
    port map (
            O => \N__41430\,
            I => \N__41421\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__41427\,
            I => \N__41417\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__41424\,
            I => \N__41414\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__41421\,
            I => \N__41411\
        );

    \I__9017\ : CEMux
    port map (
            O => \N__41420\,
            I => \N__41408\
        );

    \I__9016\ : Span4Mux_h
    port map (
            O => \N__41417\,
            I => \N__41405\
        );

    \I__9015\ : Span4Mux_h
    port map (
            O => \N__41414\,
            I => \N__41402\
        );

    \I__9014\ : Span4Mux_v
    port map (
            O => \N__41411\,
            I => \N__41399\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__41408\,
            I => \N__41396\
        );

    \I__9012\ : Span4Mux_v
    port map (
            O => \N__41405\,
            I => \N__41393\
        );

    \I__9011\ : Span4Mux_h
    port map (
            O => \N__41402\,
            I => \N__41390\
        );

    \I__9010\ : Span4Mux_h
    port map (
            O => \N__41399\,
            I => \N__41385\
        );

    \I__9009\ : Span4Mux_v
    port map (
            O => \N__41396\,
            I => \N__41385\
        );

    \I__9008\ : Odrv4
    port map (
            O => \N__41393\,
            I => \delay_measurement_inst.delay_hc_timer.N_164_i\
        );

    \I__9007\ : Odrv4
    port map (
            O => \N__41390\,
            I => \delay_measurement_inst.delay_hc_timer.N_164_i\
        );

    \I__9006\ : Odrv4
    port map (
            O => \N__41385\,
            I => \delay_measurement_inst.delay_hc_timer.N_164_i\
        );

    \I__9005\ : CascadeMux
    port map (
            O => \N__41378\,
            I => \N__41375\
        );

    \I__9004\ : InMux
    port map (
            O => \N__41375\,
            I => \N__41372\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__41372\,
            I => \N__41369\
        );

    \I__9002\ : Span4Mux_v
    port map (
            O => \N__41369\,
            I => \N__41366\
        );

    \I__9001\ : Odrv4
    port map (
            O => \N__41366\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\
        );

    \I__9000\ : InMux
    port map (
            O => \N__41363\,
            I => \N__41360\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__41360\,
            I => \N__41357\
        );

    \I__8998\ : Span4Mux_h
    port map (
            O => \N__41357\,
            I => \N__41354\
        );

    \I__8997\ : Odrv4
    port map (
            O => \N__41354\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__8996\ : CascadeMux
    port map (
            O => \N__41351\,
            I => \N__41348\
        );

    \I__8995\ : InMux
    port map (
            O => \N__41348\,
            I => \N__41345\
        );

    \I__8994\ : LocalMux
    port map (
            O => \N__41345\,
            I => \N__41342\
        );

    \I__8993\ : Odrv12
    port map (
            O => \N__41342\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\
        );

    \I__8992\ : InMux
    port map (
            O => \N__41339\,
            I => \N__41335\
        );

    \I__8991\ : InMux
    port map (
            O => \N__41338\,
            I => \N__41332\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__41335\,
            I => \N__41328\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__41332\,
            I => \N__41325\
        );

    \I__8988\ : InMux
    port map (
            O => \N__41331\,
            I => \N__41322\
        );

    \I__8987\ : Odrv4
    port map (
            O => \N__41328\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__8986\ : Odrv12
    port map (
            O => \N__41325\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__41322\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__8984\ : CascadeMux
    port map (
            O => \N__41315\,
            I => \N__41312\
        );

    \I__8983\ : InMux
    port map (
            O => \N__41312\,
            I => \N__41309\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__41309\,
            I => \N__41306\
        );

    \I__8981\ : Span4Mux_h
    port map (
            O => \N__41306\,
            I => \N__41303\
        );

    \I__8980\ : Odrv4
    port map (
            O => \N__41303\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\
        );

    \I__8979\ : CascadeMux
    port map (
            O => \N__41300\,
            I => \N__41297\
        );

    \I__8978\ : InMux
    port map (
            O => \N__41297\,
            I => \N__41294\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__41294\,
            I => \N__41291\
        );

    \I__8976\ : Span4Mux_h
    port map (
            O => \N__41291\,
            I => \N__41288\
        );

    \I__8975\ : Odrv4
    port map (
            O => \N__41288\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\
        );

    \I__8974\ : InMux
    port map (
            O => \N__41285\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__8973\ : InMux
    port map (
            O => \N__41282\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__8972\ : InMux
    port map (
            O => \N__41279\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__8971\ : InMux
    port map (
            O => \N__41276\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__8970\ : InMux
    port map (
            O => \N__41273\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__8969\ : InMux
    port map (
            O => \N__41270\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__8968\ : InMux
    port map (
            O => \N__41267\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__8967\ : InMux
    port map (
            O => \N__41264\,
            I => \bfn_17_13_0_\
        );

    \I__8966\ : InMux
    port map (
            O => \N__41261\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__8965\ : InMux
    port map (
            O => \N__41258\,
            I => \bfn_17_11_0_\
        );

    \I__8964\ : InMux
    port map (
            O => \N__41255\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__8963\ : InMux
    port map (
            O => \N__41252\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__8962\ : InMux
    port map (
            O => \N__41249\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__8961\ : InMux
    port map (
            O => \N__41246\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__8960\ : InMux
    port map (
            O => \N__41243\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__8959\ : InMux
    port map (
            O => \N__41240\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__8958\ : InMux
    port map (
            O => \N__41237\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__8957\ : InMux
    port map (
            O => \N__41234\,
            I => \bfn_17_12_0_\
        );

    \I__8956\ : CascadeMux
    port map (
            O => \N__41231\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13_cascade_\
        );

    \I__8955\ : InMux
    port map (
            O => \N__41228\,
            I => \N__41225\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__41225\,
            I => \N__41222\
        );

    \I__8953\ : Span4Mux_h
    port map (
            O => \N__41222\,
            I => \N__41219\
        );

    \I__8952\ : Odrv4
    port map (
            O => \N__41219\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__8951\ : InMux
    port map (
            O => \N__41216\,
            I => \bfn_17_10_0_\
        );

    \I__8950\ : InMux
    port map (
            O => \N__41213\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__8949\ : InMux
    port map (
            O => \N__41210\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__8948\ : InMux
    port map (
            O => \N__41207\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__8947\ : InMux
    port map (
            O => \N__41204\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__8946\ : InMux
    port map (
            O => \N__41201\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__8945\ : InMux
    port map (
            O => \N__41198\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__8944\ : InMux
    port map (
            O => \N__41195\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__8943\ : CascadeMux
    port map (
            O => \N__41192\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\
        );

    \I__8942\ : InMux
    port map (
            O => \N__41189\,
            I => \N__41186\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__41186\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\
        );

    \I__8940\ : InMux
    port map (
            O => \N__41183\,
            I => \N__41180\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__41180\,
            I => \N__41177\
        );

    \I__8938\ : Odrv4
    port map (
            O => \N__41177\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\
        );

    \I__8937\ : InMux
    port map (
            O => \N__41174\,
            I => \N__41171\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__41171\,
            I => \N__41167\
        );

    \I__8935\ : InMux
    port map (
            O => \N__41170\,
            I => \N__41163\
        );

    \I__8934\ : Span4Mux_v
    port map (
            O => \N__41167\,
            I => \N__41160\
        );

    \I__8933\ : InMux
    port map (
            O => \N__41166\,
            I => \N__41157\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__41163\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__8931\ : Odrv4
    port map (
            O => \N__41160\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__41157\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__8929\ : CascadeMux
    port map (
            O => \N__41150\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18_cascade_\
        );

    \I__8928\ : InMux
    port map (
            O => \N__41147\,
            I => \N__41144\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__41144\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\
        );

    \I__8926\ : CascadeMux
    port map (
            O => \N__41141\,
            I => \N__41138\
        );

    \I__8925\ : InMux
    port map (
            O => \N__41138\,
            I => \N__41135\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__41135\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\
        );

    \I__8923\ : InMux
    port map (
            O => \N__41132\,
            I => \N__41129\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__41129\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\
        );

    \I__8921\ : InMux
    port map (
            O => \N__41126\,
            I => \N__41123\
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__41123\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\
        );

    \I__8919\ : InMux
    port map (
            O => \N__41120\,
            I => \N__41116\
        );

    \I__8918\ : InMux
    port map (
            O => \N__41119\,
            I => \N__41113\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__41116\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__41113\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__8915\ : InMux
    port map (
            O => \N__41108\,
            I => \N__41105\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__41105\,
            I => \N__41102\
        );

    \I__8913\ : Span4Mux_h
    port map (
            O => \N__41102\,
            I => \N__41099\
        );

    \I__8912\ : Odrv4
    port map (
            O => \N__41099\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__8911\ : InMux
    port map (
            O => \N__41096\,
            I => \N__41093\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__41093\,
            I => \N__41090\
        );

    \I__8909\ : Span4Mux_v
    port map (
            O => \N__41090\,
            I => \N__41086\
        );

    \I__8908\ : InMux
    port map (
            O => \N__41089\,
            I => \N__41083\
        );

    \I__8907\ : Odrv4
    port map (
            O => \N__41086\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__41083\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__8905\ : CascadeMux
    port map (
            O => \N__41078\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\
        );

    \I__8904\ : InMux
    port map (
            O => \N__41075\,
            I => \N__41072\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__41072\,
            I => \N__41069\
        );

    \I__8902\ : Span4Mux_v
    port map (
            O => \N__41069\,
            I => \N__41066\
        );

    \I__8901\ : Odrv4
    port map (
            O => \N__41066\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__8900\ : InMux
    port map (
            O => \N__41063\,
            I => \N__41060\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__41060\,
            I => \N__41056\
        );

    \I__8898\ : InMux
    port map (
            O => \N__41059\,
            I => \N__41052\
        );

    \I__8897\ : Span4Mux_v
    port map (
            O => \N__41056\,
            I => \N__41049\
        );

    \I__8896\ : InMux
    port map (
            O => \N__41055\,
            I => \N__41046\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__41052\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__8894\ : Odrv4
    port map (
            O => \N__41049\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__41046\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__8892\ : InMux
    port map (
            O => \N__41039\,
            I => \N__41036\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__41036\,
            I => \N__41033\
        );

    \I__8890\ : Span4Mux_h
    port map (
            O => \N__41033\,
            I => \N__41030\
        );

    \I__8889\ : Odrv4
    port map (
            O => \N__41030\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__8888\ : CascadeMux
    port map (
            O => \N__41027\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\
        );

    \I__8887\ : InMux
    port map (
            O => \N__41024\,
            I => \N__41021\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__41021\,
            I => \N__41018\
        );

    \I__8885\ : Span4Mux_h
    port map (
            O => \N__41018\,
            I => \N__41015\
        );

    \I__8884\ : Odrv4
    port map (
            O => \N__41015\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\
        );

    \I__8883\ : CascadeMux
    port map (
            O => \N__41012\,
            I => \N__41009\
        );

    \I__8882\ : InMux
    port map (
            O => \N__41009\,
            I => \N__41005\
        );

    \I__8881\ : InMux
    port map (
            O => \N__41008\,
            I => \N__41002\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__41005\,
            I => \N__40998\
        );

    \I__8879\ : LocalMux
    port map (
            O => \N__41002\,
            I => \N__40995\
        );

    \I__8878\ : InMux
    port map (
            O => \N__41001\,
            I => \N__40992\
        );

    \I__8877\ : Odrv4
    port map (
            O => \N__40998\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__8876\ : Odrv12
    port map (
            O => \N__40995\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__40992\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__8874\ : CascadeMux
    port map (
            O => \N__40985\,
            I => \N__40982\
        );

    \I__8873\ : InMux
    port map (
            O => \N__40982\,
            I => \N__40979\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__40979\,
            I => \N__40976\
        );

    \I__8871\ : Odrv12
    port map (
            O => \N__40976\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt16\
        );

    \I__8870\ : InMux
    port map (
            O => \N__40973\,
            I => \N__40969\
        );

    \I__8869\ : InMux
    port map (
            O => \N__40972\,
            I => \N__40966\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__40969\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__40966\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__8866\ : InMux
    port map (
            O => \N__40961\,
            I => \N__40957\
        );

    \I__8865\ : InMux
    port map (
            O => \N__40960\,
            I => \N__40954\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__40957\,
            I => \N__40948\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__40954\,
            I => \N__40948\
        );

    \I__8862\ : InMux
    port map (
            O => \N__40953\,
            I => \N__40945\
        );

    \I__8861\ : Span4Mux_h
    port map (
            O => \N__40948\,
            I => \N__40942\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__40945\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__8859\ : Odrv4
    port map (
            O => \N__40942\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__8858\ : CascadeMux
    port map (
            O => \N__40937\,
            I => \N__40933\
        );

    \I__8857\ : InMux
    port map (
            O => \N__40936\,
            I => \N__40928\
        );

    \I__8856\ : InMux
    port map (
            O => \N__40933\,
            I => \N__40928\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__40928\,
            I => \N__40924\
        );

    \I__8854\ : InMux
    port map (
            O => \N__40927\,
            I => \N__40921\
        );

    \I__8853\ : Span4Mux_h
    port map (
            O => \N__40924\,
            I => \N__40918\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__40921\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__8851\ : Odrv4
    port map (
            O => \N__40918\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__8850\ : InMux
    port map (
            O => \N__40913\,
            I => \N__40910\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__40910\,
            I => \N__40907\
        );

    \I__8848\ : Span4Mux_h
    port map (
            O => \N__40907\,
            I => \N__40904\
        );

    \I__8847\ : Odrv4
    port map (
            O => \N__40904\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\
        );

    \I__8846\ : InMux
    port map (
            O => \N__40901\,
            I => \N__40898\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__40898\,
            I => \N__40895\
        );

    \I__8844\ : Span4Mux_v
    port map (
            O => \N__40895\,
            I => \N__40891\
        );

    \I__8843\ : InMux
    port map (
            O => \N__40894\,
            I => \N__40888\
        );

    \I__8842\ : Odrv4
    port map (
            O => \N__40891\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__40888\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__8840\ : CascadeMux
    port map (
            O => \N__40883\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\
        );

    \I__8839\ : CascadeMux
    port map (
            O => \N__40880\,
            I => \N__40877\
        );

    \I__8838\ : InMux
    port map (
            O => \N__40877\,
            I => \N__40871\
        );

    \I__8837\ : InMux
    port map (
            O => \N__40876\,
            I => \N__40871\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__40871\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__8835\ : InMux
    port map (
            O => \N__40868\,
            I => \N__40865\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__40865\,
            I => \N__40861\
        );

    \I__8833\ : InMux
    port map (
            O => \N__40864\,
            I => \N__40857\
        );

    \I__8832\ : Span4Mux_v
    port map (
            O => \N__40861\,
            I => \N__40854\
        );

    \I__8831\ : InMux
    port map (
            O => \N__40860\,
            I => \N__40851\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__40857\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__8829\ : Odrv4
    port map (
            O => \N__40854\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__40851\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__8827\ : InMux
    port map (
            O => \N__40844\,
            I => \N__40840\
        );

    \I__8826\ : InMux
    port map (
            O => \N__40843\,
            I => \N__40837\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__40840\,
            I => \N__40831\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__40837\,
            I => \N__40831\
        );

    \I__8823\ : InMux
    port map (
            O => \N__40836\,
            I => \N__40828\
        );

    \I__8822\ : Span4Mux_v
    port map (
            O => \N__40831\,
            I => \N__40825\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__40828\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__8820\ : Odrv4
    port map (
            O => \N__40825\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__8819\ : InMux
    port map (
            O => \N__40820\,
            I => \N__40817\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__40817\,
            I => \N__40814\
        );

    \I__8817\ : Span4Mux_v
    port map (
            O => \N__40814\,
            I => \N__40811\
        );

    \I__8816\ : Odrv4
    port map (
            O => \N__40811\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__8815\ : InMux
    port map (
            O => \N__40808\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__8814\ : InMux
    port map (
            O => \N__40805\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__8813\ : InMux
    port map (
            O => \N__40802\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__8812\ : InMux
    port map (
            O => \N__40799\,
            I => \bfn_16_20_0_\
        );

    \I__8811\ : InMux
    port map (
            O => \N__40796\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__8810\ : InMux
    port map (
            O => \N__40793\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__8809\ : InMux
    port map (
            O => \N__40790\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__8808\ : InMux
    port map (
            O => \N__40787\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__8807\ : InMux
    port map (
            O => \N__40784\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__8806\ : InMux
    port map (
            O => \N__40781\,
            I => \N__40778\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__40778\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__8804\ : InMux
    port map (
            O => \N__40775\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__8803\ : InMux
    port map (
            O => \N__40772\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__8802\ : InMux
    port map (
            O => \N__40769\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__8801\ : InMux
    port map (
            O => \N__40766\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__8800\ : InMux
    port map (
            O => \N__40763\,
            I => \bfn_16_19_0_\
        );

    \I__8799\ : InMux
    port map (
            O => \N__40760\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__8798\ : InMux
    port map (
            O => \N__40757\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__8797\ : InMux
    port map (
            O => \N__40754\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__8796\ : InMux
    port map (
            O => \N__40751\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__8795\ : InMux
    port map (
            O => \N__40748\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__8794\ : InMux
    port map (
            O => \N__40745\,
            I => \N__40742\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__40742\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__8792\ : InMux
    port map (
            O => \N__40739\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__8791\ : CascadeMux
    port map (
            O => \N__40736\,
            I => \N__40733\
        );

    \I__8790\ : InMux
    port map (
            O => \N__40733\,
            I => \N__40729\
        );

    \I__8789\ : InMux
    port map (
            O => \N__40732\,
            I => \N__40725\
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__40729\,
            I => \N__40722\
        );

    \I__8787\ : InMux
    port map (
            O => \N__40728\,
            I => \N__40719\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__40725\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__8785\ : Odrv12
    port map (
            O => \N__40722\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__40719\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__8783\ : InMux
    port map (
            O => \N__40712\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__8782\ : CascadeMux
    port map (
            O => \N__40709\,
            I => \N__40705\
        );

    \I__8781\ : InMux
    port map (
            O => \N__40708\,
            I => \N__40702\
        );

    \I__8780\ : InMux
    port map (
            O => \N__40705\,
            I => \N__40699\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__40702\,
            I => \N__40696\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__40699\,
            I => \N__40692\
        );

    \I__8777\ : Span4Mux_h
    port map (
            O => \N__40696\,
            I => \N__40689\
        );

    \I__8776\ : InMux
    port map (
            O => \N__40695\,
            I => \N__40686\
        );

    \I__8775\ : Odrv12
    port map (
            O => \N__40692\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__8774\ : Odrv4
    port map (
            O => \N__40689\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__40686\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__8772\ : InMux
    port map (
            O => \N__40679\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__8771\ : InMux
    port map (
            O => \N__40676\,
            I => \N__40673\
        );

    \I__8770\ : LocalMux
    port map (
            O => \N__40673\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__8769\ : InMux
    port map (
            O => \N__40670\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__8768\ : CascadeMux
    port map (
            O => \N__40667\,
            I => \N__40663\
        );

    \I__8767\ : InMux
    port map (
            O => \N__40666\,
            I => \N__40655\
        );

    \I__8766\ : InMux
    port map (
            O => \N__40663\,
            I => \N__40655\
        );

    \I__8765\ : InMux
    port map (
            O => \N__40662\,
            I => \N__40655\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__40655\,
            I => \N__40652\
        );

    \I__8763\ : Odrv4
    port map (
            O => \N__40652\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__8762\ : InMux
    port map (
            O => \N__40649\,
            I => \bfn_16_18_0_\
        );

    \I__8761\ : InMux
    port map (
            O => \N__40646\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__8760\ : InMux
    port map (
            O => \N__40643\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__8759\ : InMux
    port map (
            O => \N__40640\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__8758\ : InMux
    port map (
            O => \N__40637\,
            I => \N__40634\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__40634\,
            I => \N__40631\
        );

    \I__8756\ : Odrv4
    port map (
            O => \N__40631\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__8755\ : InMux
    port map (
            O => \N__40628\,
            I => \N__40619\
        );

    \I__8754\ : InMux
    port map (
            O => \N__40627\,
            I => \N__40619\
        );

    \I__8753\ : InMux
    port map (
            O => \N__40626\,
            I => \N__40619\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__40619\,
            I => \N__40616\
        );

    \I__8751\ : Odrv4
    port map (
            O => \N__40616\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__8750\ : InMux
    port map (
            O => \N__40613\,
            I => \N__40610\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__40610\,
            I => \N__40606\
        );

    \I__8748\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40603\
        );

    \I__8747\ : Span4Mux_h
    port map (
            O => \N__40606\,
            I => \N__40599\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__40603\,
            I => \N__40596\
        );

    \I__8745\ : InMux
    port map (
            O => \N__40602\,
            I => \N__40593\
        );

    \I__8744\ : Odrv4
    port map (
            O => \N__40599\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__8743\ : Odrv12
    port map (
            O => \N__40596\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__40593\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__8741\ : InMux
    port map (
            O => \N__40586\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__8740\ : InMux
    port map (
            O => \N__40583\,
            I => \N__40577\
        );

    \I__8739\ : InMux
    port map (
            O => \N__40582\,
            I => \N__40577\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__40577\,
            I => \N__40574\
        );

    \I__8737\ : Span4Mux_h
    port map (
            O => \N__40574\,
            I => \N__40570\
        );

    \I__8736\ : InMux
    port map (
            O => \N__40573\,
            I => \N__40567\
        );

    \I__8735\ : Odrv4
    port map (
            O => \N__40570\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__40567\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__8733\ : InMux
    port map (
            O => \N__40562\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__8732\ : InMux
    port map (
            O => \N__40559\,
            I => \N__40556\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__40556\,
            I => \N__40553\
        );

    \I__8730\ : Span4Mux_h
    port map (
            O => \N__40553\,
            I => \N__40550\
        );

    \I__8729\ : Odrv4
    port map (
            O => \N__40550\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\
        );

    \I__8728\ : InMux
    port map (
            O => \N__40547\,
            I => \N__40544\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__40544\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\
        );

    \I__8726\ : InMux
    port map (
            O => \N__40541\,
            I => \N__40538\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__40538\,
            I => \N__40535\
        );

    \I__8724\ : Span4Mux_h
    port map (
            O => \N__40535\,
            I => \N__40532\
        );

    \I__8723\ : Odrv4
    port map (
            O => \N__40532\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__8722\ : CascadeMux
    port map (
            O => \N__40529\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__8721\ : InMux
    port map (
            O => \N__40526\,
            I => \N__40523\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__40523\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\
        );

    \I__8719\ : InMux
    port map (
            O => \N__40520\,
            I => \N__40517\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__40517\,
            I => \N__40514\
        );

    \I__8717\ : Odrv4
    port map (
            O => \N__40514\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\
        );

    \I__8716\ : InMux
    port map (
            O => \N__40511\,
            I => \N__40508\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__40508\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\
        );

    \I__8714\ : CascadeMux
    port map (
            O => \N__40505\,
            I => \N__40502\
        );

    \I__8713\ : InMux
    port map (
            O => \N__40502\,
            I => \N__40499\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__40499\,
            I => \N__40496\
        );

    \I__8711\ : Span4Mux_h
    port map (
            O => \N__40496\,
            I => \N__40493\
        );

    \I__8710\ : Odrv4
    port map (
            O => \N__40493\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__8709\ : InMux
    port map (
            O => \N__40490\,
            I => \N__40483\
        );

    \I__8708\ : InMux
    port map (
            O => \N__40489\,
            I => \N__40483\
        );

    \I__8707\ : CascadeMux
    port map (
            O => \N__40488\,
            I => \N__40480\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__40483\,
            I => \N__40477\
        );

    \I__8705\ : InMux
    port map (
            O => \N__40480\,
            I => \N__40474\
        );

    \I__8704\ : Span4Mux_v
    port map (
            O => \N__40477\,
            I => \N__40470\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__40474\,
            I => \N__40467\
        );

    \I__8702\ : InMux
    port map (
            O => \N__40473\,
            I => \N__40464\
        );

    \I__8701\ : Odrv4
    port map (
            O => \N__40470\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__8700\ : Odrv4
    port map (
            O => \N__40467\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__40464\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__8698\ : InMux
    port map (
            O => \N__40457\,
            I => \N__40454\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__40454\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__8696\ : CascadeMux
    port map (
            O => \N__40451\,
            I => \N__40447\
        );

    \I__8695\ : InMux
    port map (
            O => \N__40450\,
            I => \N__40440\
        );

    \I__8694\ : InMux
    port map (
            O => \N__40447\,
            I => \N__40440\
        );

    \I__8693\ : InMux
    port map (
            O => \N__40446\,
            I => \N__40435\
        );

    \I__8692\ : InMux
    port map (
            O => \N__40445\,
            I => \N__40435\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__40440\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__40435\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8689\ : InMux
    port map (
            O => \N__40430\,
            I => \N__40427\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__40427\,
            I => \N__40424\
        );

    \I__8687\ : Odrv4
    port map (
            O => \N__40424\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__8686\ : InMux
    port map (
            O => \N__40421\,
            I => \N__40418\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__40418\,
            I => \N__40414\
        );

    \I__8684\ : InMux
    port map (
            O => \N__40417\,
            I => \N__40411\
        );

    \I__8683\ : Odrv12
    port map (
            O => \N__40414\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__40411\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__8681\ : InMux
    port map (
            O => \N__40406\,
            I => \N__40400\
        );

    \I__8680\ : InMux
    port map (
            O => \N__40405\,
            I => \N__40400\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__40400\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\
        );

    \I__8678\ : InMux
    port map (
            O => \N__40397\,
            I => \N__40394\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__40394\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__8676\ : InMux
    port map (
            O => \N__40391\,
            I => \N__40388\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__40388\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__8674\ : InMux
    port map (
            O => \N__40385\,
            I => \N__40382\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__40382\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__8672\ : InMux
    port map (
            O => \N__40379\,
            I => \N__40376\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__40376\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__8670\ : CascadeMux
    port map (
            O => \N__40373\,
            I => \N__40370\
        );

    \I__8669\ : InMux
    port map (
            O => \N__40370\,
            I => \N__40367\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__40367\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\
        );

    \I__8667\ : InMux
    port map (
            O => \N__40364\,
            I => \N__40361\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__40361\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\
        );

    \I__8665\ : InMux
    port map (
            O => \N__40358\,
            I => \N__40355\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__40355\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\
        );

    \I__8663\ : CascadeMux
    port map (
            O => \N__40352\,
            I => \N__40349\
        );

    \I__8662\ : InMux
    port map (
            O => \N__40349\,
            I => \N__40346\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__40346\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\
        );

    \I__8660\ : CascadeMux
    port map (
            O => \N__40343\,
            I => \N__40340\
        );

    \I__8659\ : InMux
    port map (
            O => \N__40340\,
            I => \N__40337\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__40337\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt20\
        );

    \I__8657\ : InMux
    port map (
            O => \N__40334\,
            I => \N__40328\
        );

    \I__8656\ : InMux
    port map (
            O => \N__40333\,
            I => \N__40328\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__40328\,
            I => \N__40324\
        );

    \I__8654\ : InMux
    port map (
            O => \N__40327\,
            I => \N__40321\
        );

    \I__8653\ : Span4Mux_h
    port map (
            O => \N__40324\,
            I => \N__40318\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__40321\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__8651\ : Odrv4
    port map (
            O => \N__40318\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__8650\ : CascadeMux
    port map (
            O => \N__40313\,
            I => \N__40310\
        );

    \I__8649\ : InMux
    port map (
            O => \N__40310\,
            I => \N__40304\
        );

    \I__8648\ : InMux
    port map (
            O => \N__40309\,
            I => \N__40304\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__40304\,
            I => \N__40300\
        );

    \I__8646\ : InMux
    port map (
            O => \N__40303\,
            I => \N__40297\
        );

    \I__8645\ : Span4Mux_h
    port map (
            O => \N__40300\,
            I => \N__40294\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__40297\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__8643\ : Odrv4
    port map (
            O => \N__40294\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__8642\ : InMux
    port map (
            O => \N__40289\,
            I => \N__40286\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__40286\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\
        );

    \I__8640\ : InMux
    port map (
            O => \N__40283\,
            I => \N__40280\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__40280\,
            I => \N__40277\
        );

    \I__8638\ : Span4Mux_v
    port map (
            O => \N__40277\,
            I => \N__40273\
        );

    \I__8637\ : InMux
    port map (
            O => \N__40276\,
            I => \N__40270\
        );

    \I__8636\ : Odrv4
    port map (
            O => \N__40273\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__40270\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__8634\ : InMux
    port map (
            O => \N__40265\,
            I => \N__40259\
        );

    \I__8633\ : InMux
    port map (
            O => \N__40264\,
            I => \N__40259\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__40259\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\
        );

    \I__8631\ : InMux
    port map (
            O => \N__40256\,
            I => \N__40253\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__40253\,
            I => \N__40250\
        );

    \I__8629\ : Span4Mux_v
    port map (
            O => \N__40250\,
            I => \N__40245\
        );

    \I__8628\ : InMux
    port map (
            O => \N__40249\,
            I => \N__40242\
        );

    \I__8627\ : InMux
    port map (
            O => \N__40248\,
            I => \N__40239\
        );

    \I__8626\ : Span4Mux_h
    port map (
            O => \N__40245\,
            I => \N__40234\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__40242\,
            I => \N__40234\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__40239\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__8623\ : Odrv4
    port map (
            O => \N__40234\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__8622\ : CascadeMux
    port map (
            O => \N__40229\,
            I => \N__40226\
        );

    \I__8621\ : InMux
    port map (
            O => \N__40226\,
            I => \N__40220\
        );

    \I__8620\ : InMux
    port map (
            O => \N__40225\,
            I => \N__40220\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__40220\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\
        );

    \I__8618\ : InMux
    port map (
            O => \N__40217\,
            I => \N__40212\
        );

    \I__8617\ : InMux
    port map (
            O => \N__40216\,
            I => \N__40209\
        );

    \I__8616\ : InMux
    port map (
            O => \N__40215\,
            I => \N__40206\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__40212\,
            I => \N__40203\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__40209\,
            I => \N__40200\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__40206\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__8612\ : Odrv12
    port map (
            O => \N__40203\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__8611\ : Odrv4
    port map (
            O => \N__40200\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__8610\ : CascadeMux
    port map (
            O => \N__40193\,
            I => \N__40190\
        );

    \I__8609\ : InMux
    port map (
            O => \N__40190\,
            I => \N__40187\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__40187\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__8607\ : InMux
    port map (
            O => \N__40184\,
            I => \N__40181\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__40181\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__8605\ : CascadeMux
    port map (
            O => \N__40178\,
            I => \N__40175\
        );

    \I__8604\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40172\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__40172\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt22\
        );

    \I__8602\ : CascadeMux
    port map (
            O => \N__40169\,
            I => \N__40165\
        );

    \I__8601\ : InMux
    port map (
            O => \N__40168\,
            I => \N__40159\
        );

    \I__8600\ : InMux
    port map (
            O => \N__40165\,
            I => \N__40159\
        );

    \I__8599\ : InMux
    port map (
            O => \N__40164\,
            I => \N__40156\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__40159\,
            I => \N__40153\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__40156\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__8596\ : Odrv4
    port map (
            O => \N__40153\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__8595\ : CascadeMux
    port map (
            O => \N__40148\,
            I => \N__40143\
        );

    \I__8594\ : InMux
    port map (
            O => \N__40147\,
            I => \N__40140\
        );

    \I__8593\ : InMux
    port map (
            O => \N__40146\,
            I => \N__40135\
        );

    \I__8592\ : InMux
    port map (
            O => \N__40143\,
            I => \N__40135\
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__40140\,
            I => \N__40130\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__40135\,
            I => \N__40130\
        );

    \I__8589\ : Odrv4
    port map (
            O => \N__40130\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__8588\ : InMux
    port map (
            O => \N__40127\,
            I => \N__40124\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__40124\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\
        );

    \I__8586\ : InMux
    port map (
            O => \N__40121\,
            I => \N__40118\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__40118\,
            I => \N__40115\
        );

    \I__8584\ : Span4Mux_v
    port map (
            O => \N__40115\,
            I => \N__40111\
        );

    \I__8583\ : InMux
    port map (
            O => \N__40114\,
            I => \N__40108\
        );

    \I__8582\ : Odrv4
    port map (
            O => \N__40111\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__40108\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__8580\ : InMux
    port map (
            O => \N__40103\,
            I => \N__40097\
        );

    \I__8579\ : InMux
    port map (
            O => \N__40102\,
            I => \N__40097\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__40097\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\
        );

    \I__8577\ : CascadeMux
    port map (
            O => \N__40094\,
            I => \N__40091\
        );

    \I__8576\ : InMux
    port map (
            O => \N__40091\,
            I => \N__40088\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__40088\,
            I => \N__40085\
        );

    \I__8574\ : Odrv4
    port map (
            O => \N__40085\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__8573\ : InMux
    port map (
            O => \N__40082\,
            I => \N__40079\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__40079\,
            I => \N__40076\
        );

    \I__8571\ : Span4Mux_h
    port map (
            O => \N__40076\,
            I => \N__40073\
        );

    \I__8570\ : Odrv4
    port map (
            O => \N__40073\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt26\
        );

    \I__8569\ : InMux
    port map (
            O => \N__40070\,
            I => \N__40064\
        );

    \I__8568\ : InMux
    port map (
            O => \N__40069\,
            I => \N__40064\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__40064\,
            I => \N__40060\
        );

    \I__8566\ : InMux
    port map (
            O => \N__40063\,
            I => \N__40057\
        );

    \I__8565\ : Span4Mux_h
    port map (
            O => \N__40060\,
            I => \N__40054\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__40057\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__8563\ : Odrv4
    port map (
            O => \N__40054\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__8562\ : CascadeMux
    port map (
            O => \N__40049\,
            I => \N__40046\
        );

    \I__8561\ : InMux
    port map (
            O => \N__40046\,
            I => \N__40040\
        );

    \I__8560\ : InMux
    port map (
            O => \N__40045\,
            I => \N__40040\
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__40040\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__8558\ : CascadeMux
    port map (
            O => \N__40037\,
            I => \N__40033\
        );

    \I__8557\ : InMux
    port map (
            O => \N__40036\,
            I => \N__40028\
        );

    \I__8556\ : InMux
    port map (
            O => \N__40033\,
            I => \N__40028\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__40028\,
            I => \N__40024\
        );

    \I__8554\ : InMux
    port map (
            O => \N__40027\,
            I => \N__40021\
        );

    \I__8553\ : Span4Mux_h
    port map (
            O => \N__40024\,
            I => \N__40018\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__40021\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__8551\ : Odrv4
    port map (
            O => \N__40018\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__8550\ : CascadeMux
    port map (
            O => \N__40013\,
            I => \N__40010\
        );

    \I__8549\ : InMux
    port map (
            O => \N__40010\,
            I => \N__40007\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__40007\,
            I => \N__40004\
        );

    \I__8547\ : Odrv4
    port map (
            O => \N__40004\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\
        );

    \I__8546\ : InMux
    port map (
            O => \N__40001\,
            I => \N__39997\
        );

    \I__8545\ : InMux
    port map (
            O => \N__40000\,
            I => \N__39993\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__39997\,
            I => \N__39990\
        );

    \I__8543\ : InMux
    port map (
            O => \N__39996\,
            I => \N__39987\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__39993\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__8541\ : Odrv12
    port map (
            O => \N__39990\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__39987\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__8539\ : InMux
    port map (
            O => \N__39980\,
            I => \N__39974\
        );

    \I__8538\ : InMux
    port map (
            O => \N__39979\,
            I => \N__39974\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__39974\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__8536\ : InMux
    port map (
            O => \N__39971\,
            I => \N__39968\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__39968\,
            I => \N__39964\
        );

    \I__8534\ : InMux
    port map (
            O => \N__39967\,
            I => \N__39961\
        );

    \I__8533\ : Odrv12
    port map (
            O => \N__39964\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__39961\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__8531\ : CascadeMux
    port map (
            O => \N__39956\,
            I => \N__39953\
        );

    \I__8530\ : InMux
    port map (
            O => \N__39953\,
            I => \N__39950\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__39950\,
            I => \N__39947\
        );

    \I__8528\ : Odrv4
    port map (
            O => \N__39947\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\
        );

    \I__8527\ : InMux
    port map (
            O => \N__39944\,
            I => \N__39938\
        );

    \I__8526\ : InMux
    port map (
            O => \N__39943\,
            I => \N__39938\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__39938\,
            I => \N__39934\
        );

    \I__8524\ : InMux
    port map (
            O => \N__39937\,
            I => \N__39931\
        );

    \I__8523\ : Span4Mux_h
    port map (
            O => \N__39934\,
            I => \N__39928\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__39931\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__8521\ : Odrv4
    port map (
            O => \N__39928\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__8520\ : CascadeMux
    port map (
            O => \N__39923\,
            I => \N__39920\
        );

    \I__8519\ : InMux
    port map (
            O => \N__39920\,
            I => \N__39914\
        );

    \I__8518\ : InMux
    port map (
            O => \N__39919\,
            I => \N__39914\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__39914\,
            I => \N__39910\
        );

    \I__8516\ : InMux
    port map (
            O => \N__39913\,
            I => \N__39907\
        );

    \I__8515\ : Span4Mux_v
    port map (
            O => \N__39910\,
            I => \N__39904\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__39907\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__8513\ : Odrv4
    port map (
            O => \N__39904\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__8512\ : InMux
    port map (
            O => \N__39899\,
            I => \N__39893\
        );

    \I__8511\ : InMux
    port map (
            O => \N__39898\,
            I => \N__39893\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__39893\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\
        );

    \I__8509\ : InMux
    port map (
            O => \N__39890\,
            I => \N__39887\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__39887\,
            I => \N__39884\
        );

    \I__8507\ : Span4Mux_h
    port map (
            O => \N__39884\,
            I => \N__39881\
        );

    \I__8506\ : Odrv4
    port map (
            O => \N__39881\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt28\
        );

    \I__8505\ : InMux
    port map (
            O => \N__39878\,
            I => \N__39875\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__39875\,
            I => \N__39871\
        );

    \I__8503\ : InMux
    port map (
            O => \N__39874\,
            I => \N__39868\
        );

    \I__8502\ : Odrv12
    port map (
            O => \N__39871\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__39868\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__8500\ : CascadeMux
    port map (
            O => \N__39863\,
            I => \N__39860\
        );

    \I__8499\ : InMux
    port map (
            O => \N__39860\,
            I => \N__39854\
        );

    \I__8498\ : InMux
    port map (
            O => \N__39859\,
            I => \N__39854\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__39854\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\
        );

    \I__8496\ : CascadeMux
    port map (
            O => \N__39851\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\
        );

    \I__8495\ : CascadeMux
    port map (
            O => \N__39848\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30_cascade_\
        );

    \I__8494\ : InMux
    port map (
            O => \N__39845\,
            I => \N__39839\
        );

    \I__8493\ : InMux
    port map (
            O => \N__39844\,
            I => \N__39839\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__39839\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\
        );

    \I__8491\ : InMux
    port map (
            O => \N__39836\,
            I => \N__39831\
        );

    \I__8490\ : InMux
    port map (
            O => \N__39835\,
            I => \N__39826\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39834\,
            I => \N__39826\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__39831\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__39826\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__8486\ : InMux
    port map (
            O => \N__39821\,
            I => \N__39816\
        );

    \I__8485\ : InMux
    port map (
            O => \N__39820\,
            I => \N__39811\
        );

    \I__8484\ : InMux
    port map (
            O => \N__39819\,
            I => \N__39811\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__39816\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__39811\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__8481\ : InMux
    port map (
            O => \N__39806\,
            I => \N__39803\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__39803\,
            I => \N__39800\
        );

    \I__8479\ : Span4Mux_h
    port map (
            O => \N__39800\,
            I => \N__39797\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__39797\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\
        );

    \I__8477\ : InMux
    port map (
            O => \N__39794\,
            I => \N__39791\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__39791\,
            I => \N__39788\
        );

    \I__8475\ : Span4Mux_h
    port map (
            O => \N__39788\,
            I => \N__39785\
        );

    \I__8474\ : Odrv4
    port map (
            O => \N__39785\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__8473\ : InMux
    port map (
            O => \N__39782\,
            I => \N__39779\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__39779\,
            I => \N__39776\
        );

    \I__8471\ : Odrv4
    port map (
            O => \N__39776\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt16\
        );

    \I__8470\ : InMux
    port map (
            O => \N__39773\,
            I => \N__39767\
        );

    \I__8469\ : InMux
    port map (
            O => \N__39772\,
            I => \N__39767\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__39767\,
            I => \N__39763\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39766\,
            I => \N__39760\
        );

    \I__8466\ : Span4Mux_h
    port map (
            O => \N__39763\,
            I => \N__39757\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__39760\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__8464\ : Odrv4
    port map (
            O => \N__39757\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__8463\ : CascadeMux
    port map (
            O => \N__39752\,
            I => \N__39748\
        );

    \I__8462\ : InMux
    port map (
            O => \N__39751\,
            I => \N__39743\
        );

    \I__8461\ : InMux
    port map (
            O => \N__39748\,
            I => \N__39743\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__39743\,
            I => \N__39739\
        );

    \I__8459\ : InMux
    port map (
            O => \N__39742\,
            I => \N__39736\
        );

    \I__8458\ : Span4Mux_h
    port map (
            O => \N__39739\,
            I => \N__39733\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__39736\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__8456\ : Odrv4
    port map (
            O => \N__39733\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__8455\ : CascadeMux
    port map (
            O => \N__39728\,
            I => \N__39725\
        );

    \I__8454\ : InMux
    port map (
            O => \N__39725\,
            I => \N__39722\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__39722\,
            I => \N__39719\
        );

    \I__8452\ : Span4Mux_h
    port map (
            O => \N__39719\,
            I => \N__39716\
        );

    \I__8451\ : Odrv4
    port map (
            O => \N__39716\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\
        );

    \I__8450\ : InMux
    port map (
            O => \N__39713\,
            I => \N__39707\
        );

    \I__8449\ : InMux
    port map (
            O => \N__39712\,
            I => \N__39707\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__39707\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__8447\ : CascadeMux
    port map (
            O => \N__39704\,
            I => \N__39701\
        );

    \I__8446\ : InMux
    port map (
            O => \N__39701\,
            I => \N__39695\
        );

    \I__8445\ : InMux
    port map (
            O => \N__39700\,
            I => \N__39695\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__39695\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__8443\ : CascadeMux
    port map (
            O => \N__39692\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\
        );

    \I__8442\ : InMux
    port map (
            O => \N__39689\,
            I => \N__39683\
        );

    \I__8441\ : InMux
    port map (
            O => \N__39688\,
            I => \N__39683\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__39683\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\
        );

    \I__8439\ : InMux
    port map (
            O => \N__39680\,
            I => \N__39677\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__39677\,
            I => \N__39674\
        );

    \I__8437\ : Span4Mux_v
    port map (
            O => \N__39674\,
            I => \N__39671\
        );

    \I__8436\ : Odrv4
    port map (
            O => \N__39671\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt22\
        );

    \I__8435\ : InMux
    port map (
            O => \N__39668\,
            I => \N__39663\
        );

    \I__8434\ : InMux
    port map (
            O => \N__39667\,
            I => \N__39658\
        );

    \I__8433\ : InMux
    port map (
            O => \N__39666\,
            I => \N__39658\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__39663\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__39658\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__8430\ : CascadeMux
    port map (
            O => \N__39653\,
            I => \N__39649\
        );

    \I__8429\ : InMux
    port map (
            O => \N__39652\,
            I => \N__39645\
        );

    \I__8428\ : InMux
    port map (
            O => \N__39649\,
            I => \N__39640\
        );

    \I__8427\ : InMux
    port map (
            O => \N__39648\,
            I => \N__39640\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__39645\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__39640\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__8424\ : CascadeMux
    port map (
            O => \N__39635\,
            I => \N__39632\
        );

    \I__8423\ : InMux
    port map (
            O => \N__39632\,
            I => \N__39629\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__39629\,
            I => \N__39626\
        );

    \I__8421\ : Span4Mux_v
    port map (
            O => \N__39626\,
            I => \N__39623\
        );

    \I__8420\ : Span4Mux_h
    port map (
            O => \N__39623\,
            I => \N__39620\
        );

    \I__8419\ : Odrv4
    port map (
            O => \N__39620\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\
        );

    \I__8418\ : CascadeMux
    port map (
            O => \N__39617\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\
        );

    \I__8417\ : CascadeMux
    port map (
            O => \N__39614\,
            I => \N__39611\
        );

    \I__8416\ : InMux
    port map (
            O => \N__39611\,
            I => \N__39605\
        );

    \I__8415\ : InMux
    port map (
            O => \N__39610\,
            I => \N__39605\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__39605\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\
        );

    \I__8413\ : CascadeMux
    port map (
            O => \N__39602\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\
        );

    \I__8412\ : InMux
    port map (
            O => \N__39599\,
            I => \N__39593\
        );

    \I__8411\ : InMux
    port map (
            O => \N__39598\,
            I => \N__39593\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__39593\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\
        );

    \I__8409\ : CascadeMux
    port map (
            O => \N__39590\,
            I => \N__39587\
        );

    \I__8408\ : InMux
    port map (
            O => \N__39587\,
            I => \N__39584\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__39584\,
            I => \N__39581\
        );

    \I__8406\ : Span4Mux_h
    port map (
            O => \N__39581\,
            I => \N__39578\
        );

    \I__8405\ : Odrv4
    port map (
            O => \N__39578\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__8404\ : InMux
    port map (
            O => \N__39575\,
            I => \N__39572\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__39572\,
            I => \N__39568\
        );

    \I__8402\ : InMux
    port map (
            O => \N__39571\,
            I => \N__39564\
        );

    \I__8401\ : Span4Mux_v
    port map (
            O => \N__39568\,
            I => \N__39561\
        );

    \I__8400\ : InMux
    port map (
            O => \N__39567\,
            I => \N__39558\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__39564\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__8398\ : Odrv4
    port map (
            O => \N__39561\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__39558\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__8396\ : InMux
    port map (
            O => \N__39551\,
            I => \N__39546\
        );

    \I__8395\ : InMux
    port map (
            O => \N__39550\,
            I => \N__39543\
        );

    \I__8394\ : CascadeMux
    port map (
            O => \N__39549\,
            I => \N__39538\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__39546\,
            I => \N__39535\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__39543\,
            I => \N__39532\
        );

    \I__8391\ : InMux
    port map (
            O => \N__39542\,
            I => \N__39527\
        );

    \I__8390\ : InMux
    port map (
            O => \N__39541\,
            I => \N__39527\
        );

    \I__8389\ : InMux
    port map (
            O => \N__39538\,
            I => \N__39524\
        );

    \I__8388\ : Span4Mux_h
    port map (
            O => \N__39535\,
            I => \N__39521\
        );

    \I__8387\ : Span4Mux_h
    port map (
            O => \N__39532\,
            I => \N__39518\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__39527\,
            I => \N__39515\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__39524\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__8384\ : Odrv4
    port map (
            O => \N__39521\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__8383\ : Odrv4
    port map (
            O => \N__39518\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__8382\ : Odrv12
    port map (
            O => \N__39515\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__8381\ : InMux
    port map (
            O => \N__39506\,
            I => \N__39501\
        );

    \I__8380\ : InMux
    port map (
            O => \N__39505\,
            I => \N__39498\
        );

    \I__8379\ : InMux
    port map (
            O => \N__39504\,
            I => \N__39495\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__39501\,
            I => \N__39492\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__39498\,
            I => \N__39489\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__39495\,
            I => \N__39486\
        );

    \I__8375\ : Span4Mux_h
    port map (
            O => \N__39492\,
            I => \N__39483\
        );

    \I__8374\ : Odrv4
    port map (
            O => \N__39489\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__8373\ : Odrv4
    port map (
            O => \N__39486\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__8372\ : Odrv4
    port map (
            O => \N__39483\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__8371\ : InMux
    port map (
            O => \N__39476\,
            I => \N__39473\
        );

    \I__8370\ : LocalMux
    port map (
            O => \N__39473\,
            I => \N__39470\
        );

    \I__8369\ : Span4Mux_h
    port map (
            O => \N__39470\,
            I => \N__39466\
        );

    \I__8368\ : InMux
    port map (
            O => \N__39469\,
            I => \N__39463\
        );

    \I__8367\ : Odrv4
    port map (
            O => \N__39466\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__39463\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__8365\ : CascadeMux
    port map (
            O => \N__39458\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__8364\ : CascadeMux
    port map (
            O => \N__39455\,
            I => \N__39452\
        );

    \I__8363\ : InMux
    port map (
            O => \N__39452\,
            I => \N__39447\
        );

    \I__8362\ : InMux
    port map (
            O => \N__39451\,
            I => \N__39442\
        );

    \I__8361\ : InMux
    port map (
            O => \N__39450\,
            I => \N__39442\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__39447\,
            I => \N__39439\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__39442\,
            I => \N__39434\
        );

    \I__8358\ : Span4Mux_h
    port map (
            O => \N__39439\,
            I => \N__39431\
        );

    \I__8357\ : InMux
    port map (
            O => \N__39438\,
            I => \N__39426\
        );

    \I__8356\ : InMux
    port map (
            O => \N__39437\,
            I => \N__39426\
        );

    \I__8355\ : Odrv4
    port map (
            O => \N__39434\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__8354\ : Odrv4
    port map (
            O => \N__39431\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__39426\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__8352\ : InMux
    port map (
            O => \N__39419\,
            I => \N__39416\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__39416\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\
        );

    \I__8350\ : CascadeMux
    port map (
            O => \N__39413\,
            I => \N__39410\
        );

    \I__8349\ : InMux
    port map (
            O => \N__39410\,
            I => \N__39407\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__39407\,
            I => \N__39404\
        );

    \I__8347\ : Span4Mux_h
    port map (
            O => \N__39404\,
            I => \N__39401\
        );

    \I__8346\ : Odrv4
    port map (
            O => \N__39401\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt28\
        );

    \I__8345\ : InMux
    port map (
            O => \N__39398\,
            I => \N__39391\
        );

    \I__8344\ : InMux
    port map (
            O => \N__39397\,
            I => \N__39391\
        );

    \I__8343\ : InMux
    port map (
            O => \N__39396\,
            I => \N__39388\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__39391\,
            I => \N__39385\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__39388\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__8340\ : Odrv4
    port map (
            O => \N__39385\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__8339\ : CascadeMux
    port map (
            O => \N__39380\,
            I => \N__39377\
        );

    \I__8338\ : InMux
    port map (
            O => \N__39377\,
            I => \N__39371\
        );

    \I__8337\ : InMux
    port map (
            O => \N__39376\,
            I => \N__39371\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__39371\,
            I => \N__39367\
        );

    \I__8335\ : InMux
    port map (
            O => \N__39370\,
            I => \N__39364\
        );

    \I__8334\ : Span4Mux_v
    port map (
            O => \N__39367\,
            I => \N__39361\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__39364\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__8332\ : Odrv4
    port map (
            O => \N__39361\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__8331\ : InMux
    port map (
            O => \N__39356\,
            I => \N__39353\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__39353\,
            I => \N__39350\
        );

    \I__8329\ : Odrv4
    port map (
            O => \N__39350\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\
        );

    \I__8328\ : CascadeMux
    port map (
            O => \N__39347\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\
        );

    \I__8327\ : CascadeMux
    port map (
            O => \N__39344\,
            I => \N__39341\
        );

    \I__8326\ : InMux
    port map (
            O => \N__39341\,
            I => \N__39335\
        );

    \I__8325\ : InMux
    port map (
            O => \N__39340\,
            I => \N__39335\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__39335\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\
        );

    \I__8323\ : InMux
    port map (
            O => \N__39332\,
            I => \N__39329\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__39329\,
            I => \N__39326\
        );

    \I__8321\ : Odrv4
    port map (
            O => \N__39326\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__8320\ : InMux
    port map (
            O => \N__39323\,
            I => \N__39320\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__39320\,
            I => \N__39317\
        );

    \I__8318\ : Odrv12
    port map (
            O => \N__39317\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__8317\ : CascadeMux
    port map (
            O => \N__39314\,
            I => \N__39311\
        );

    \I__8316\ : InMux
    port map (
            O => \N__39311\,
            I => \N__39308\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__39308\,
            I => \N__39305\
        );

    \I__8314\ : Span4Mux_v
    port map (
            O => \N__39305\,
            I => \N__39302\
        );

    \I__8313\ : Odrv4
    port map (
            O => \N__39302\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__8312\ : InMux
    port map (
            O => \N__39299\,
            I => \N__39296\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__39296\,
            I => \N__39293\
        );

    \I__8310\ : Span4Mux_h
    port map (
            O => \N__39293\,
            I => \N__39289\
        );

    \I__8309\ : InMux
    port map (
            O => \N__39292\,
            I => \N__39285\
        );

    \I__8308\ : Span4Mux_v
    port map (
            O => \N__39289\,
            I => \N__39282\
        );

    \I__8307\ : InMux
    port map (
            O => \N__39288\,
            I => \N__39279\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__39285\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__8305\ : Odrv4
    port map (
            O => \N__39282\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__39279\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__8303\ : InMux
    port map (
            O => \N__39272\,
            I => \N__39268\
        );

    \I__8302\ : InMux
    port map (
            O => \N__39271\,
            I => \N__39265\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__39268\,
            I => \N__39262\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__39265\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__8299\ : Odrv4
    port map (
            O => \N__39262\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__8298\ : CascadeMux
    port map (
            O => \N__39257\,
            I => \N__39252\
        );

    \I__8297\ : InMux
    port map (
            O => \N__39256\,
            I => \N__39246\
        );

    \I__8296\ : InMux
    port map (
            O => \N__39255\,
            I => \N__39246\
        );

    \I__8295\ : InMux
    port map (
            O => \N__39252\,
            I => \N__39241\
        );

    \I__8294\ : InMux
    port map (
            O => \N__39251\,
            I => \N__39241\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__39246\,
            I => \N__39238\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__39241\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8291\ : Odrv12
    port map (
            O => \N__39238\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8290\ : InMux
    port map (
            O => \N__39233\,
            I => \N__39229\
        );

    \I__8289\ : InMux
    port map (
            O => \N__39232\,
            I => \N__39225\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__39229\,
            I => \N__39222\
        );

    \I__8287\ : InMux
    port map (
            O => \N__39228\,
            I => \N__39219\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__39225\,
            I => \N__39214\
        );

    \I__8285\ : Span4Mux_v
    port map (
            O => \N__39222\,
            I => \N__39214\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__39219\,
            I => \N__39211\
        );

    \I__8283\ : Odrv4
    port map (
            O => \N__39214\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__8282\ : Odrv12
    port map (
            O => \N__39211\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__8281\ : CascadeMux
    port map (
            O => \N__39206\,
            I => \N__39203\
        );

    \I__8280\ : InMux
    port map (
            O => \N__39203\,
            I => \N__39200\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__39200\,
            I => \N__39197\
        );

    \I__8278\ : Odrv4
    port map (
            O => \N__39197\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30\
        );

    \I__8277\ : CascadeMux
    port map (
            O => \N__39194\,
            I => \N__39191\
        );

    \I__8276\ : InMux
    port map (
            O => \N__39191\,
            I => \N__39188\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__39188\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__8274\ : InMux
    port map (
            O => \N__39185\,
            I => \N__39182\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__39182\,
            I => \N__39179\
        );

    \I__8272\ : Odrv12
    port map (
            O => \N__39179\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\
        );

    \I__8271\ : CascadeMux
    port map (
            O => \N__39176\,
            I => \N__39173\
        );

    \I__8270\ : InMux
    port map (
            O => \N__39173\,
            I => \N__39170\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__39170\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__8268\ : InMux
    port map (
            O => \N__39167\,
            I => \N__39164\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__39164\,
            I => \N__39161\
        );

    \I__8266\ : Odrv4
    port map (
            O => \N__39161\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__8265\ : InMux
    port map (
            O => \N__39158\,
            I => \N__39155\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__39155\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__8263\ : InMux
    port map (
            O => \N__39152\,
            I => \N__39149\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__39149\,
            I => \N__39146\
        );

    \I__8261\ : Odrv4
    port map (
            O => \N__39146\,
            I => \current_shift_inst.control_input_axb_23\
        );

    \I__8260\ : CascadeMux
    port map (
            O => \N__39143\,
            I => \N__39140\
        );

    \I__8259\ : InMux
    port map (
            O => \N__39140\,
            I => \N__39137\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__39137\,
            I => \N__39134\
        );

    \I__8257\ : Odrv4
    port map (
            O => \N__39134\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__8256\ : CascadeMux
    port map (
            O => \N__39131\,
            I => \N__39128\
        );

    \I__8255\ : InMux
    port map (
            O => \N__39128\,
            I => \N__39125\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__39125\,
            I => \N__39122\
        );

    \I__8253\ : Span4Mux_v
    port map (
            O => \N__39122\,
            I => \N__39119\
        );

    \I__8252\ : Odrv4
    port map (
            O => \N__39119\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\
        );

    \I__8251\ : CascadeMux
    port map (
            O => \N__39116\,
            I => \N__39113\
        );

    \I__8250\ : InMux
    port map (
            O => \N__39113\,
            I => \N__39110\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__39110\,
            I => \N__39107\
        );

    \I__8248\ : Span4Mux_h
    port map (
            O => \N__39107\,
            I => \N__39104\
        );

    \I__8247\ : Odrv4
    port map (
            O => \N__39104\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__8246\ : CascadeMux
    port map (
            O => \N__39101\,
            I => \N__39098\
        );

    \I__8245\ : InMux
    port map (
            O => \N__39098\,
            I => \N__39095\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__39095\,
            I => \N__39092\
        );

    \I__8243\ : Odrv12
    port map (
            O => \N__39092\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__8242\ : CascadeMux
    port map (
            O => \N__39089\,
            I => \N__39086\
        );

    \I__8241\ : InMux
    port map (
            O => \N__39086\,
            I => \N__39083\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__39083\,
            I => \N__39080\
        );

    \I__8239\ : Span4Mux_v
    port map (
            O => \N__39080\,
            I => \N__39077\
        );

    \I__8238\ : Odrv4
    port map (
            O => \N__39077\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\
        );

    \I__8237\ : InMux
    port map (
            O => \N__39074\,
            I => \N__39071\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__39071\,
            I => \current_shift_inst.un38_control_input_0_s0_16\
        );

    \I__8235\ : InMux
    port map (
            O => \N__39068\,
            I => \N__39065\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__39065\,
            I => \N__39062\
        );

    \I__8233\ : Odrv12
    port map (
            O => \N__39062\,
            I => \current_shift_inst.un38_control_input_0_s1_16\
        );

    \I__8232\ : InMux
    port map (
            O => \N__39059\,
            I => \N__39056\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__39056\,
            I => \N__39053\
        );

    \I__8230\ : Odrv4
    port map (
            O => \N__39053\,
            I => \current_shift_inst.control_input_axb_13\
        );

    \I__8229\ : InMux
    port map (
            O => \N__39050\,
            I => \N__39047\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__39047\,
            I => \current_shift_inst.un38_control_input_0_s0_17\
        );

    \I__8227\ : InMux
    port map (
            O => \N__39044\,
            I => \N__39041\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__39041\,
            I => \N__39038\
        );

    \I__8225\ : Span4Mux_v
    port map (
            O => \N__39038\,
            I => \N__39035\
        );

    \I__8224\ : Odrv4
    port map (
            O => \N__39035\,
            I => \current_shift_inst.un38_control_input_0_s1_17\
        );

    \I__8223\ : InMux
    port map (
            O => \N__39032\,
            I => \N__39029\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__39029\,
            I => \N__39026\
        );

    \I__8221\ : Odrv4
    port map (
            O => \N__39026\,
            I => \current_shift_inst.control_input_axb_14\
        );

    \I__8220\ : InMux
    port map (
            O => \N__39023\,
            I => \N__39020\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__39020\,
            I => \N__39017\
        );

    \I__8218\ : Odrv4
    port map (
            O => \N__39017\,
            I => \current_shift_inst.un38_control_input_0_s1_18\
        );

    \I__8217\ : InMux
    port map (
            O => \N__39014\,
            I => \N__39011\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__39011\,
            I => \current_shift_inst.un38_control_input_0_s0_18\
        );

    \I__8215\ : InMux
    port map (
            O => \N__39008\,
            I => \N__39005\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__39005\,
            I => \N__39002\
        );

    \I__8213\ : Odrv4
    port map (
            O => \N__39002\,
            I => \current_shift_inst.control_input_axb_15\
        );

    \I__8212\ : InMux
    port map (
            O => \N__38999\,
            I => \N__38996\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__38996\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\
        );

    \I__8210\ : InMux
    port map (
            O => \N__38993\,
            I => \N__38990\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__38990\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__8208\ : CascadeMux
    port map (
            O => \N__38987\,
            I => \N__38984\
        );

    \I__8207\ : InMux
    port map (
            O => \N__38984\,
            I => \N__38981\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__38981\,
            I => \N__38978\
        );

    \I__8205\ : Odrv12
    port map (
            O => \N__38978\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__8204\ : InMux
    port map (
            O => \N__38975\,
            I => \N__38972\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__38972\,
            I => \N__38969\
        );

    \I__8202\ : Odrv4
    port map (
            O => \N__38969\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__8201\ : CascadeMux
    port map (
            O => \N__38966\,
            I => \N__38963\
        );

    \I__8200\ : InMux
    port map (
            O => \N__38963\,
            I => \N__38960\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__38960\,
            I => \N__38957\
        );

    \I__8198\ : Odrv4
    port map (
            O => \N__38957\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__8197\ : InMux
    port map (
            O => \N__38954\,
            I => \N__38951\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__38951\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__8195\ : CascadeMux
    port map (
            O => \N__38948\,
            I => \N__38945\
        );

    \I__8194\ : InMux
    port map (
            O => \N__38945\,
            I => \N__38942\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__38942\,
            I => \N__38939\
        );

    \I__8192\ : Span4Mux_v
    port map (
            O => \N__38939\,
            I => \N__38936\
        );

    \I__8191\ : Odrv4
    port map (
            O => \N__38936\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__38933\,
            I => \N__38930\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38930\,
            I => \N__38927\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__38927\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\
        );

    \I__8187\ : CascadeMux
    port map (
            O => \N__38924\,
            I => \N__38921\
        );

    \I__8186\ : InMux
    port map (
            O => \N__38921\,
            I => \N__38918\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__38918\,
            I => \N__38915\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__38915\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\
        );

    \I__8183\ : InMux
    port map (
            O => \N__38912\,
            I => \N__38909\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__38909\,
            I => \N__38906\
        );

    \I__8181\ : Odrv12
    port map (
            O => \N__38906\,
            I => \current_shift_inst.un38_control_input_0_s1_15\
        );

    \I__8180\ : InMux
    port map (
            O => \N__38903\,
            I => \N__38900\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__38900\,
            I => \N__38897\
        );

    \I__8178\ : Odrv4
    port map (
            O => \N__38897\,
            I => \current_shift_inst.un38_control_input_0_s0_15\
        );

    \I__8177\ : InMux
    port map (
            O => \N__38894\,
            I => \N__38891\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__38891\,
            I => \N__38888\
        );

    \I__8175\ : Odrv12
    port map (
            O => \N__38888\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__8174\ : InMux
    port map (
            O => \N__38885\,
            I => \N__38882\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__38882\,
            I => \N__38879\
        );

    \I__8172\ : Odrv12
    port map (
            O => \N__38879\,
            I => \current_shift_inst.un38_control_input_0_s1_14\
        );

    \I__8171\ : InMux
    port map (
            O => \N__38876\,
            I => \N__38873\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__38873\,
            I => \N__38870\
        );

    \I__8169\ : Odrv4
    port map (
            O => \N__38870\,
            I => \current_shift_inst.un38_control_input_0_s0_14\
        );

    \I__8168\ : InMux
    port map (
            O => \N__38867\,
            I => \N__38864\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__38864\,
            I => \N__38861\
        );

    \I__8166\ : Odrv12
    port map (
            O => \N__38861\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__8165\ : InMux
    port map (
            O => \N__38858\,
            I => \N__38855\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__38855\,
            I => \N__38852\
        );

    \I__8163\ : Odrv4
    port map (
            O => \N__38852\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38849\,
            I => \N__38846\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__38846\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__8160\ : InMux
    port map (
            O => \N__38843\,
            I => \N__38840\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__38840\,
            I => \N__38837\
        );

    \I__8158\ : Span4Mux_v
    port map (
            O => \N__38837\,
            I => \N__38834\
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__38834\,
            I => \current_shift_inst.control_input_axb_24\
        );

    \I__8156\ : InMux
    port map (
            O => \N__38831\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__8155\ : InMux
    port map (
            O => \N__38828\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__8154\ : InMux
    port map (
            O => \N__38825\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__8153\ : InMux
    port map (
            O => \N__38822\,
            I => \N__38819\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__38819\,
            I => \N__38816\
        );

    \I__8151\ : Span4Mux_h
    port map (
            O => \N__38816\,
            I => \N__38813\
        );

    \I__8150\ : Span4Mux_v
    port map (
            O => \N__38813\,
            I => \N__38810\
        );

    \I__8149\ : Odrv4
    port map (
            O => \N__38810\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__8148\ : InMux
    port map (
            O => \N__38807\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__8147\ : InMux
    port map (
            O => \N__38804\,
            I => \N__38801\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__38801\,
            I => \N__38798\
        );

    \I__8145\ : Span4Mux_v
    port map (
            O => \N__38798\,
            I => \N__38795\
        );

    \I__8144\ : Sp12to4
    port map (
            O => \N__38795\,
            I => \N__38792\
        );

    \I__8143\ : Odrv12
    port map (
            O => \N__38792\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__8142\ : InMux
    port map (
            O => \N__38789\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38786\,
            I => \N__38783\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__38783\,
            I => \N__38780\
        );

    \I__8139\ : Span4Mux_h
    port map (
            O => \N__38780\,
            I => \N__38777\
        );

    \I__8138\ : Odrv4
    port map (
            O => \N__38777\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__8137\ : InMux
    port map (
            O => \N__38774\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__8136\ : InMux
    port map (
            O => \N__38771\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__8135\ : InMux
    port map (
            O => \N__38768\,
            I => \N__38765\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__38765\,
            I => \N__38762\
        );

    \I__8133\ : Span4Mux_v
    port map (
            O => \N__38762\,
            I => \N__38759\
        );

    \I__8132\ : Sp12to4
    port map (
            O => \N__38759\,
            I => \N__38756\
        );

    \I__8131\ : Odrv12
    port map (
            O => \N__38756\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38753\,
            I => \N__38750\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__38750\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38747\,
            I => \N__38744\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__38744\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\
        );

    \I__8126\ : InMux
    port map (
            O => \N__38741\,
            I => \current_shift_inst.un38_control_input_cry_16_s1\
        );

    \I__8125\ : InMux
    port map (
            O => \N__38738\,
            I => \current_shift_inst.un38_control_input_cry_17_s1\
        );

    \I__8124\ : CascadeMux
    port map (
            O => \N__38735\,
            I => \N__38732\
        );

    \I__8123\ : InMux
    port map (
            O => \N__38732\,
            I => \N__38729\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__38729\,
            I => \N__38726\
        );

    \I__8121\ : Span4Mux_h
    port map (
            O => \N__38726\,
            I => \N__38723\
        );

    \I__8120\ : Odrv4
    port map (
            O => \N__38723\,
            I => \current_shift_inst.un38_control_input_0_s1_19\
        );

    \I__8119\ : InMux
    port map (
            O => \N__38720\,
            I => \current_shift_inst.un38_control_input_cry_18_s1\
        );

    \I__8118\ : CascadeMux
    port map (
            O => \N__38717\,
            I => \N__38714\
        );

    \I__8117\ : InMux
    port map (
            O => \N__38714\,
            I => \N__38711\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__38711\,
            I => \N__38708\
        );

    \I__8115\ : Span4Mux_v
    port map (
            O => \N__38708\,
            I => \N__38705\
        );

    \I__8114\ : Odrv4
    port map (
            O => \N__38705\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__8113\ : InMux
    port map (
            O => \N__38702\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__8112\ : InMux
    port map (
            O => \N__38699\,
            I => \N__38696\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__38696\,
            I => \N__38693\
        );

    \I__8110\ : Span4Mux_v
    port map (
            O => \N__38693\,
            I => \N__38690\
        );

    \I__8109\ : Odrv4
    port map (
            O => \N__38690\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__8108\ : InMux
    port map (
            O => \N__38687\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__8107\ : InMux
    port map (
            O => \N__38684\,
            I => \N__38681\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__38681\,
            I => \N__38678\
        );

    \I__8105\ : Span4Mux_v
    port map (
            O => \N__38678\,
            I => \N__38675\
        );

    \I__8104\ : Odrv4
    port map (
            O => \N__38675\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__8103\ : InMux
    port map (
            O => \N__38672\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__8102\ : CascadeMux
    port map (
            O => \N__38669\,
            I => \N__38666\
        );

    \I__8101\ : InMux
    port map (
            O => \N__38666\,
            I => \N__38663\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__38663\,
            I => \N__38660\
        );

    \I__8099\ : Span4Mux_v
    port map (
            O => \N__38660\,
            I => \N__38657\
        );

    \I__8098\ : Odrv4
    port map (
            O => \N__38657\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__8097\ : InMux
    port map (
            O => \N__38654\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__8096\ : InMux
    port map (
            O => \N__38651\,
            I => \N__38648\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__38648\,
            I => \N__38645\
        );

    \I__8094\ : Span4Mux_v
    port map (
            O => \N__38645\,
            I => \N__38642\
        );

    \I__8093\ : Odrv4
    port map (
            O => \N__38642\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__8092\ : InMux
    port map (
            O => \N__38639\,
            I => \bfn_15_16_0_\
        );

    \I__8091\ : InMux
    port map (
            O => \N__38636\,
            I => \N__38633\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__38633\,
            I => \N__38630\
        );

    \I__8089\ : Span4Mux_v
    port map (
            O => \N__38630\,
            I => \N__38627\
        );

    \I__8088\ : Odrv4
    port map (
            O => \N__38627\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__8087\ : InMux
    port map (
            O => \N__38624\,
            I => \N__38621\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__38621\,
            I => \N__38618\
        );

    \I__8085\ : Span4Mux_v
    port map (
            O => \N__38618\,
            I => \N__38615\
        );

    \I__8084\ : Odrv4
    port map (
            O => \N__38615\,
            I => \current_shift_inst.un38_control_input_0_s1_8\
        );

    \I__8083\ : InMux
    port map (
            O => \N__38612\,
            I => \bfn_15_14_0_\
        );

    \I__8082\ : InMux
    port map (
            O => \N__38609\,
            I => \N__38606\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__38606\,
            I => \N__38603\
        );

    \I__8080\ : Span4Mux_v
    port map (
            O => \N__38603\,
            I => \N__38600\
        );

    \I__8079\ : Odrv4
    port map (
            O => \N__38600\,
            I => \current_shift_inst.un38_control_input_0_s1_9\
        );

    \I__8078\ : InMux
    port map (
            O => \N__38597\,
            I => \current_shift_inst.un38_control_input_cry_8_s1\
        );

    \I__8077\ : InMux
    port map (
            O => \N__38594\,
            I => \N__38591\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__38591\,
            I => \N__38588\
        );

    \I__8075\ : Span4Mux_v
    port map (
            O => \N__38588\,
            I => \N__38585\
        );

    \I__8074\ : Odrv4
    port map (
            O => \N__38585\,
            I => \current_shift_inst.un38_control_input_0_s1_10\
        );

    \I__8073\ : InMux
    port map (
            O => \N__38582\,
            I => \current_shift_inst.un38_control_input_cry_9_s1\
        );

    \I__8072\ : InMux
    port map (
            O => \N__38579\,
            I => \N__38576\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__38576\,
            I => \N__38573\
        );

    \I__8070\ : Span4Mux_v
    port map (
            O => \N__38573\,
            I => \N__38570\
        );

    \I__8069\ : Odrv4
    port map (
            O => \N__38570\,
            I => \current_shift_inst.un38_control_input_0_s1_11\
        );

    \I__8068\ : InMux
    port map (
            O => \N__38567\,
            I => \current_shift_inst.un38_control_input_cry_10_s1\
        );

    \I__8067\ : InMux
    port map (
            O => \N__38564\,
            I => \N__38561\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__38561\,
            I => \N__38558\
        );

    \I__8065\ : Span12Mux_h
    port map (
            O => \N__38558\,
            I => \N__38555\
        );

    \I__8064\ : Odrv12
    port map (
            O => \N__38555\,
            I => \current_shift_inst.un38_control_input_0_s1_12\
        );

    \I__8063\ : InMux
    port map (
            O => \N__38552\,
            I => \current_shift_inst.un38_control_input_cry_11_s1\
        );

    \I__8062\ : InMux
    port map (
            O => \N__38549\,
            I => \N__38546\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__38546\,
            I => \N__38543\
        );

    \I__8060\ : Span4Mux_v
    port map (
            O => \N__38543\,
            I => \N__38540\
        );

    \I__8059\ : Odrv4
    port map (
            O => \N__38540\,
            I => \current_shift_inst.un38_control_input_0_s1_13\
        );

    \I__8058\ : InMux
    port map (
            O => \N__38537\,
            I => \current_shift_inst.un38_control_input_cry_12_s1\
        );

    \I__8057\ : InMux
    port map (
            O => \N__38534\,
            I => \current_shift_inst.un38_control_input_cry_13_s1\
        );

    \I__8056\ : InMux
    port map (
            O => \N__38531\,
            I => \current_shift_inst.un38_control_input_cry_14_s1\
        );

    \I__8055\ : InMux
    port map (
            O => \N__38528\,
            I => \bfn_15_15_0_\
        );

    \I__8054\ : CascadeMux
    port map (
            O => \N__38525\,
            I => \N__38522\
        );

    \I__8053\ : InMux
    port map (
            O => \N__38522\,
            I => \N__38519\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__38519\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\
        );

    \I__8051\ : InMux
    port map (
            O => \N__38516\,
            I => \N__38513\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__38513\,
            I => \N__38510\
        );

    \I__8049\ : Span4Mux_v
    port map (
            O => \N__38510\,
            I => \N__38507\
        );

    \I__8048\ : Span4Mux_h
    port map (
            O => \N__38507\,
            I => \N__38504\
        );

    \I__8047\ : Odrv4
    port map (
            O => \N__38504\,
            I => \current_shift_inst.un38_control_input_0_s1_3\
        );

    \I__8046\ : InMux
    port map (
            O => \N__38501\,
            I => \current_shift_inst.un38_control_input_cry_2_s1\
        );

    \I__8045\ : InMux
    port map (
            O => \N__38498\,
            I => \N__38495\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__38495\,
            I => \N__38492\
        );

    \I__8043\ : Span4Mux_v
    port map (
            O => \N__38492\,
            I => \N__38489\
        );

    \I__8042\ : Span4Mux_v
    port map (
            O => \N__38489\,
            I => \N__38486\
        );

    \I__8041\ : Odrv4
    port map (
            O => \N__38486\,
            I => \current_shift_inst.un38_control_input_0_s1_4\
        );

    \I__8040\ : InMux
    port map (
            O => \N__38483\,
            I => \current_shift_inst.un38_control_input_cry_3_s1\
        );

    \I__8039\ : CascadeMux
    port map (
            O => \N__38480\,
            I => \N__38477\
        );

    \I__8038\ : InMux
    port map (
            O => \N__38477\,
            I => \N__38474\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__38474\,
            I => \N__38471\
        );

    \I__8036\ : Span12Mux_h
    port map (
            O => \N__38471\,
            I => \N__38468\
        );

    \I__8035\ : Odrv12
    port map (
            O => \N__38468\,
            I => \current_shift_inst.un38_control_input_0_s1_5\
        );

    \I__8034\ : InMux
    port map (
            O => \N__38465\,
            I => \current_shift_inst.un38_control_input_cry_4_s1\
        );

    \I__8033\ : InMux
    port map (
            O => \N__38462\,
            I => \N__38459\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__38459\,
            I => \N__38456\
        );

    \I__8031\ : Span12Mux_v
    port map (
            O => \N__38456\,
            I => \N__38453\
        );

    \I__8030\ : Odrv12
    port map (
            O => \N__38453\,
            I => \current_shift_inst.un38_control_input_0_s1_6\
        );

    \I__8029\ : InMux
    port map (
            O => \N__38450\,
            I => \current_shift_inst.un38_control_input_cry_5_s1\
        );

    \I__8028\ : InMux
    port map (
            O => \N__38447\,
            I => \N__38444\
        );

    \I__8027\ : LocalMux
    port map (
            O => \N__38444\,
            I => \N__38441\
        );

    \I__8026\ : Span4Mux_h
    port map (
            O => \N__38441\,
            I => \N__38438\
        );

    \I__8025\ : Span4Mux_v
    port map (
            O => \N__38438\,
            I => \N__38435\
        );

    \I__8024\ : Odrv4
    port map (
            O => \N__38435\,
            I => \current_shift_inst.un38_control_input_0_s1_7\
        );

    \I__8023\ : InMux
    port map (
            O => \N__38432\,
            I => \current_shift_inst.un38_control_input_cry_6_s1\
        );

    \I__8022\ : InMux
    port map (
            O => \N__38429\,
            I => \N__38426\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__38426\,
            I => \N__38423\
        );

    \I__8020\ : Span4Mux_v
    port map (
            O => \N__38423\,
            I => \N__38420\
        );

    \I__8019\ : Odrv4
    port map (
            O => \N__38420\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\
        );

    \I__8018\ : CascadeMux
    port map (
            O => \N__38417\,
            I => \N__38414\
        );

    \I__8017\ : InMux
    port map (
            O => \N__38414\,
            I => \N__38411\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__38411\,
            I => \N__38408\
        );

    \I__8015\ : Span4Mux_v
    port map (
            O => \N__38408\,
            I => \N__38405\
        );

    \I__8014\ : Odrv4
    port map (
            O => \N__38405\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt18\
        );

    \I__8013\ : InMux
    port map (
            O => \N__38402\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30\
        );

    \I__8012\ : CascadeMux
    port map (
            O => \N__38399\,
            I => \N__38396\
        );

    \I__8011\ : InMux
    port map (
            O => \N__38396\,
            I => \N__38393\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__38393\,
            I => \N__38388\
        );

    \I__8009\ : InMux
    port map (
            O => \N__38392\,
            I => \N__38385\
        );

    \I__8008\ : InMux
    port map (
            O => \N__38391\,
            I => \N__38382\
        );

    \I__8007\ : Span4Mux_h
    port map (
            O => \N__38388\,
            I => \N__38379\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__38385\,
            I => \N__38376\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__38382\,
            I => \N__38373\
        );

    \I__8004\ : Span4Mux_h
    port map (
            O => \N__38379\,
            I => \N__38370\
        );

    \I__8003\ : Span4Mux_h
    port map (
            O => \N__38376\,
            I => \N__38367\
        );

    \I__8002\ : Span4Mux_v
    port map (
            O => \N__38373\,
            I => \N__38364\
        );

    \I__8001\ : Span4Mux_v
    port map (
            O => \N__38370\,
            I => \N__38361\
        );

    \I__8000\ : Span4Mux_h
    port map (
            O => \N__38367\,
            I => \N__38358\
        );

    \I__7999\ : Odrv4
    port map (
            O => \N__38364\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__7998\ : Odrv4
    port map (
            O => \N__38361\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__7997\ : Odrv4
    port map (
            O => \N__38358\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__7996\ : InMux
    port map (
            O => \N__38351\,
            I => \N__38348\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__38348\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__7994\ : InMux
    port map (
            O => \N__38345\,
            I => \N__38341\
        );

    \I__7993\ : InMux
    port map (
            O => \N__38344\,
            I => \N__38338\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__38341\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__38338\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__7990\ : CascadeMux
    port map (
            O => \N__38333\,
            I => \N__38330\
        );

    \I__7989\ : InMux
    port map (
            O => \N__38330\,
            I => \N__38327\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__38327\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__7987\ : InMux
    port map (
            O => \N__38324\,
            I => \N__38320\
        );

    \I__7986\ : InMux
    port map (
            O => \N__38323\,
            I => \N__38317\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__38320\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__38317\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__7983\ : CascadeMux
    port map (
            O => \N__38312\,
            I => \N__38309\
        );

    \I__7982\ : InMux
    port map (
            O => \N__38309\,
            I => \N__38306\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__38306\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__7980\ : InMux
    port map (
            O => \N__38303\,
            I => \N__38299\
        );

    \I__7979\ : InMux
    port map (
            O => \N__38302\,
            I => \N__38296\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__38299\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__38296\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7976\ : CascadeMux
    port map (
            O => \N__38291\,
            I => \N__38288\
        );

    \I__7975\ : InMux
    port map (
            O => \N__38288\,
            I => \N__38285\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__38285\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__7973\ : InMux
    port map (
            O => \N__38282\,
            I => \N__38278\
        );

    \I__7972\ : InMux
    port map (
            O => \N__38281\,
            I => \N__38275\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__38278\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__38275\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7969\ : CascadeMux
    port map (
            O => \N__38270\,
            I => \N__38267\
        );

    \I__7968\ : InMux
    port map (
            O => \N__38267\,
            I => \N__38264\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__38264\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__7966\ : InMux
    port map (
            O => \N__38261\,
            I => \N__38257\
        );

    \I__7965\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38254\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__38257\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__38254\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7962\ : CascadeMux
    port map (
            O => \N__38249\,
            I => \N__38246\
        );

    \I__7961\ : InMux
    port map (
            O => \N__38246\,
            I => \N__38243\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__38243\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__7959\ : InMux
    port map (
            O => \N__38240\,
            I => \N__38236\
        );

    \I__7958\ : InMux
    port map (
            O => \N__38239\,
            I => \N__38233\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__38236\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__38233\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__7955\ : CascadeMux
    port map (
            O => \N__38228\,
            I => \N__38225\
        );

    \I__7954\ : InMux
    port map (
            O => \N__38225\,
            I => \N__38222\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__38222\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__7952\ : InMux
    port map (
            O => \N__38219\,
            I => \N__38215\
        );

    \I__7951\ : InMux
    port map (
            O => \N__38218\,
            I => \N__38212\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__38215\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__38212\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7948\ : InMux
    port map (
            O => \N__38207\,
            I => \N__38204\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__38204\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__7946\ : CascadeMux
    port map (
            O => \N__38201\,
            I => \N__38198\
        );

    \I__7945\ : InMux
    port map (
            O => \N__38198\,
            I => \N__38195\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__38195\,
            I => \N__38192\
        );

    \I__7943\ : Odrv4
    port map (
            O => \N__38192\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__7942\ : InMux
    port map (
            O => \N__38189\,
            I => \N__38185\
        );

    \I__7941\ : InMux
    port map (
            O => \N__38188\,
            I => \N__38182\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__38185\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__38182\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__7938\ : InMux
    port map (
            O => \N__38177\,
            I => \N__38174\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__38174\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__7936\ : CascadeMux
    port map (
            O => \N__38171\,
            I => \N__38168\
        );

    \I__7935\ : InMux
    port map (
            O => \N__38168\,
            I => \N__38165\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__38165\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__7933\ : CascadeMux
    port map (
            O => \N__38162\,
            I => \N__38158\
        );

    \I__7932\ : InMux
    port map (
            O => \N__38161\,
            I => \N__38154\
        );

    \I__7931\ : InMux
    port map (
            O => \N__38158\,
            I => \N__38151\
        );

    \I__7930\ : InMux
    port map (
            O => \N__38157\,
            I => \N__38148\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__38154\,
            I => \N__38145\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__38151\,
            I => \N__38142\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__38148\,
            I => \N__38137\
        );

    \I__7926\ : Span4Mux_h
    port map (
            O => \N__38145\,
            I => \N__38137\
        );

    \I__7925\ : Odrv12
    port map (
            O => \N__38142\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7924\ : Odrv4
    port map (
            O => \N__38137\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7923\ : InMux
    port map (
            O => \N__38132\,
            I => \N__38129\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__38129\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__7921\ : InMux
    port map (
            O => \N__38126\,
            I => \N__38123\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__38123\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__7919\ : InMux
    port map (
            O => \N__38120\,
            I => \N__38116\
        );

    \I__7918\ : InMux
    port map (
            O => \N__38119\,
            I => \N__38113\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__38116\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__38113\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__7915\ : CascadeMux
    port map (
            O => \N__38108\,
            I => \N__38105\
        );

    \I__7914\ : InMux
    port map (
            O => \N__38105\,
            I => \N__38102\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__38102\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__7912\ : CascadeMux
    port map (
            O => \N__38099\,
            I => \N__38096\
        );

    \I__7911\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38093\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__38093\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__7909\ : InMux
    port map (
            O => \N__38090\,
            I => \N__38086\
        );

    \I__7908\ : InMux
    port map (
            O => \N__38089\,
            I => \N__38083\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__38086\,
            I => \N__38080\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__38083\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7905\ : Odrv4
    port map (
            O => \N__38080\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7904\ : InMux
    port map (
            O => \N__38075\,
            I => \N__38072\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__38072\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__7902\ : InMux
    port map (
            O => \N__38069\,
            I => \N__38065\
        );

    \I__7901\ : InMux
    port map (
            O => \N__38068\,
            I => \N__38062\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__38065\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__38062\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7898\ : InMux
    port map (
            O => \N__38057\,
            I => \N__38054\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__38054\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__7896\ : CascadeMux
    port map (
            O => \N__38051\,
            I => \N__38048\
        );

    \I__7895\ : InMux
    port map (
            O => \N__38048\,
            I => \N__38045\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__38045\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__7893\ : InMux
    port map (
            O => \N__38042\,
            I => \N__38039\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__38039\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__7891\ : InMux
    port map (
            O => \N__38036\,
            I => \N__38032\
        );

    \I__7890\ : InMux
    port map (
            O => \N__38035\,
            I => \N__38029\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__38032\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__38029\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7887\ : CascadeMux
    port map (
            O => \N__38024\,
            I => \N__38021\
        );

    \I__7886\ : InMux
    port map (
            O => \N__38021\,
            I => \N__38018\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__38018\,
            I => \N__38015\
        );

    \I__7884\ : Odrv4
    port map (
            O => \N__38015\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__7883\ : InMux
    port map (
            O => \N__38012\,
            I => \N__38008\
        );

    \I__7882\ : InMux
    port map (
            O => \N__38011\,
            I => \N__38005\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__38008\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__38005\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7879\ : InMux
    port map (
            O => \N__38000\,
            I => \N__37997\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__37997\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__7877\ : CascadeMux
    port map (
            O => \N__37994\,
            I => \N__37991\
        );

    \I__7876\ : InMux
    port map (
            O => \N__37991\,
            I => \N__37988\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__37988\,
            I => \N__37985\
        );

    \I__7874\ : Odrv4
    port map (
            O => \N__37985\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__7873\ : InMux
    port map (
            O => \N__37982\,
            I => \N__37978\
        );

    \I__7872\ : InMux
    port map (
            O => \N__37981\,
            I => \N__37975\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__37978\,
            I => \N__37972\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__37975\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__7869\ : Odrv4
    port map (
            O => \N__37972\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__7868\ : InMux
    port map (
            O => \N__37967\,
            I => \N__37964\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__37964\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__7866\ : InMux
    port map (
            O => \N__37961\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__7865\ : InMux
    port map (
            O => \N__37958\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__7864\ : InMux
    port map (
            O => \N__37955\,
            I => \N__37952\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__37952\,
            I => \N__37949\
        );

    \I__7862\ : Span4Mux_h
    port map (
            O => \N__37949\,
            I => \N__37945\
        );

    \I__7861\ : InMux
    port map (
            O => \N__37948\,
            I => \N__37942\
        );

    \I__7860\ : Odrv4
    port map (
            O => \N__37945\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__37942\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__7858\ : InMux
    port map (
            O => \N__37937\,
            I => \N__37932\
        );

    \I__7857\ : InMux
    port map (
            O => \N__37936\,
            I => \N__37929\
        );

    \I__7856\ : InMux
    port map (
            O => \N__37935\,
            I => \N__37926\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__37932\,
            I => \N__37923\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__37929\,
            I => \N__37918\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__37926\,
            I => \N__37918\
        );

    \I__7852\ : Odrv12
    port map (
            O => \N__37923\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__7851\ : Odrv4
    port map (
            O => \N__37918\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__7850\ : InMux
    port map (
            O => \N__37913\,
            I => \N__37908\
        );

    \I__7849\ : InMux
    port map (
            O => \N__37912\,
            I => \N__37905\
        );

    \I__7848\ : InMux
    port map (
            O => \N__37911\,
            I => \N__37902\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__37908\,
            I => \N__37899\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__37905\,
            I => \N__37896\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__37902\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__7844\ : Odrv4
    port map (
            O => \N__37899\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__7843\ : Odrv4
    port map (
            O => \N__37896\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__7842\ : InMux
    port map (
            O => \N__37889\,
            I => \N__37885\
        );

    \I__7841\ : InMux
    port map (
            O => \N__37888\,
            I => \N__37882\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__37885\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__37882\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__7838\ : InMux
    port map (
            O => \N__37877\,
            I => \N__37873\
        );

    \I__7837\ : InMux
    port map (
            O => \N__37876\,
            I => \N__37869\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__37873\,
            I => \N__37866\
        );

    \I__7835\ : InMux
    port map (
            O => \N__37872\,
            I => \N__37863\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__37869\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__7833\ : Odrv4
    port map (
            O => \N__37866\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__37863\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__7831\ : InMux
    port map (
            O => \N__37856\,
            I => \N__37852\
        );

    \I__7830\ : InMux
    port map (
            O => \N__37855\,
            I => \N__37848\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__37852\,
            I => \N__37845\
        );

    \I__7828\ : InMux
    port map (
            O => \N__37851\,
            I => \N__37842\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__37848\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__7826\ : Odrv4
    port map (
            O => \N__37845\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__37842\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__7824\ : InMux
    port map (
            O => \N__37835\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__7823\ : InMux
    port map (
            O => \N__37832\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__7822\ : InMux
    port map (
            O => \N__37829\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__7821\ : InMux
    port map (
            O => \N__37826\,
            I => \N__37823\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__37823\,
            I => \N__37818\
        );

    \I__7819\ : InMux
    port map (
            O => \N__37822\,
            I => \N__37815\
        );

    \I__7818\ : InMux
    port map (
            O => \N__37821\,
            I => \N__37812\
        );

    \I__7817\ : Span4Mux_h
    port map (
            O => \N__37818\,
            I => \N__37809\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__37815\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__37812\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__7814\ : Odrv4
    port map (
            O => \N__37809\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__7813\ : InMux
    port map (
            O => \N__37802\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__7812\ : InMux
    port map (
            O => \N__37799\,
            I => \N__37795\
        );

    \I__7811\ : CascadeMux
    port map (
            O => \N__37798\,
            I => \N__37791\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__37795\,
            I => \N__37788\
        );

    \I__7809\ : InMux
    port map (
            O => \N__37794\,
            I => \N__37785\
        );

    \I__7808\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37782\
        );

    \I__7807\ : Span4Mux_h
    port map (
            O => \N__37788\,
            I => \N__37779\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__37785\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__37782\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__7804\ : Odrv4
    port map (
            O => \N__37779\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37772\,
            I => \bfn_15_8_0_\
        );

    \I__7802\ : CascadeMux
    port map (
            O => \N__37769\,
            I => \N__37765\
        );

    \I__7801\ : InMux
    port map (
            O => \N__37768\,
            I => \N__37761\
        );

    \I__7800\ : InMux
    port map (
            O => \N__37765\,
            I => \N__37756\
        );

    \I__7799\ : InMux
    port map (
            O => \N__37764\,
            I => \N__37756\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__37761\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__37756\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__7796\ : InMux
    port map (
            O => \N__37751\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__7795\ : InMux
    port map (
            O => \N__37748\,
            I => \N__37743\
        );

    \I__7794\ : InMux
    port map (
            O => \N__37747\,
            I => \N__37738\
        );

    \I__7793\ : InMux
    port map (
            O => \N__37746\,
            I => \N__37738\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__37743\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__37738\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__7790\ : InMux
    port map (
            O => \N__37733\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__7789\ : InMux
    port map (
            O => \N__37730\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__7788\ : InMux
    port map (
            O => \N__37727\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__7787\ : InMux
    port map (
            O => \N__37724\,
            I => \N__37720\
        );

    \I__7786\ : InMux
    port map (
            O => \N__37723\,
            I => \N__37717\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__37720\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__37717\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7783\ : InMux
    port map (
            O => \N__37712\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__7782\ : InMux
    port map (
            O => \N__37709\,
            I => \N__37705\
        );

    \I__7781\ : InMux
    port map (
            O => \N__37708\,
            I => \N__37702\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__37705\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__37702\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__7778\ : InMux
    port map (
            O => \N__37697\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__7777\ : InMux
    port map (
            O => \N__37694\,
            I => \N__37690\
        );

    \I__7776\ : InMux
    port map (
            O => \N__37693\,
            I => \N__37687\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__37690\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__37687\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7773\ : InMux
    port map (
            O => \N__37682\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__7772\ : InMux
    port map (
            O => \N__37679\,
            I => \N__37675\
        );

    \I__7771\ : InMux
    port map (
            O => \N__37678\,
            I => \N__37672\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__37675\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__37672\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__7768\ : InMux
    port map (
            O => \N__37667\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__7767\ : InMux
    port map (
            O => \N__37664\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__7766\ : InMux
    port map (
            O => \N__37661\,
            I => \bfn_15_7_0_\
        );

    \I__7765\ : CascadeMux
    port map (
            O => \N__37658\,
            I => \N__37654\
        );

    \I__7764\ : InMux
    port map (
            O => \N__37657\,
            I => \N__37650\
        );

    \I__7763\ : InMux
    port map (
            O => \N__37654\,
            I => \N__37647\
        );

    \I__7762\ : InMux
    port map (
            O => \N__37653\,
            I => \N__37644\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__37650\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__37647\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__37644\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7758\ : InMux
    port map (
            O => \N__37637\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__7757\ : InMux
    port map (
            O => \N__37634\,
            I => \N__37629\
        );

    \I__7756\ : InMux
    port map (
            O => \N__37633\,
            I => \N__37626\
        );

    \I__7755\ : InMux
    port map (
            O => \N__37632\,
            I => \N__37623\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__37629\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__37626\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__37623\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7751\ : InMux
    port map (
            O => \N__37616\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__7750\ : CascadeMux
    port map (
            O => \N__37613\,
            I => \N__37609\
        );

    \I__7749\ : CascadeMux
    port map (
            O => \N__37612\,
            I => \N__37605\
        );

    \I__7748\ : InMux
    port map (
            O => \N__37609\,
            I => \N__37602\
        );

    \I__7747\ : InMux
    port map (
            O => \N__37608\,
            I => \N__37599\
        );

    \I__7746\ : InMux
    port map (
            O => \N__37605\,
            I => \N__37596\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__37602\,
            I => \N__37593\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__37599\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__37596\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__7742\ : Odrv4
    port map (
            O => \N__37593\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__7741\ : InMux
    port map (
            O => \N__37586\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__7740\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37579\
        );

    \I__7739\ : InMux
    port map (
            O => \N__37582\,
            I => \N__37576\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__37579\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__37576\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7736\ : InMux
    port map (
            O => \N__37571\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__7735\ : InMux
    port map (
            O => \N__37568\,
            I => \N__37564\
        );

    \I__7734\ : InMux
    port map (
            O => \N__37567\,
            I => \N__37561\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__37564\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__37561\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7731\ : InMux
    port map (
            O => \N__37556\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__7730\ : InMux
    port map (
            O => \N__37553\,
            I => \N__37549\
        );

    \I__7729\ : InMux
    port map (
            O => \N__37552\,
            I => \N__37546\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__37549\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__37546\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7726\ : InMux
    port map (
            O => \N__37541\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__7725\ : InMux
    port map (
            O => \N__37538\,
            I => \N__37534\
        );

    \I__7724\ : InMux
    port map (
            O => \N__37537\,
            I => \N__37531\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__37534\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__37531\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__7721\ : InMux
    port map (
            O => \N__37526\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__7720\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37519\
        );

    \I__7719\ : InMux
    port map (
            O => \N__37522\,
            I => \N__37516\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__37519\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__37516\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__7716\ : InMux
    port map (
            O => \N__37511\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__7715\ : InMux
    port map (
            O => \N__37508\,
            I => \N__37504\
        );

    \I__7714\ : InMux
    port map (
            O => \N__37507\,
            I => \N__37501\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__37504\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__37501\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__7711\ : InMux
    port map (
            O => \N__37496\,
            I => \bfn_15_6_0_\
        );

    \I__7710\ : InMux
    port map (
            O => \N__37493\,
            I => \N__37489\
        );

    \I__7709\ : InMux
    port map (
            O => \N__37492\,
            I => \N__37486\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__37489\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__37486\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7706\ : InMux
    port map (
            O => \N__37481\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__7705\ : InMux
    port map (
            O => \N__37478\,
            I => \N__37474\
        );

    \I__7704\ : InMux
    port map (
            O => \N__37477\,
            I => \N__37471\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__37474\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__37471\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7701\ : InMux
    port map (
            O => \N__37466\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__7700\ : InMux
    port map (
            O => \N__37463\,
            I => \N__37457\
        );

    \I__7699\ : InMux
    port map (
            O => \N__37462\,
            I => \N__37452\
        );

    \I__7698\ : InMux
    port map (
            O => \N__37461\,
            I => \N__37452\
        );

    \I__7697\ : InMux
    port map (
            O => \N__37460\,
            I => \N__37449\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__37457\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__37452\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__37449\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7693\ : InMux
    port map (
            O => \N__37442\,
            I => \N__37436\
        );

    \I__7692\ : InMux
    port map (
            O => \N__37441\,
            I => \N__37431\
        );

    \I__7691\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37431\
        );

    \I__7690\ : InMux
    port map (
            O => \N__37439\,
            I => \N__37428\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__37436\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__37431\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__37428\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7686\ : CascadeMux
    port map (
            O => \N__37421\,
            I => \N__37417\
        );

    \I__7685\ : InMux
    port map (
            O => \N__37420\,
            I => \N__37412\
        );

    \I__7684\ : InMux
    port map (
            O => \N__37417\,
            I => \N__37409\
        );

    \I__7683\ : InMux
    port map (
            O => \N__37416\,
            I => \N__37406\
        );

    \I__7682\ : InMux
    port map (
            O => \N__37415\,
            I => \N__37403\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__37412\,
            I => \N__37400\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__37409\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__37406\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__37403\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7677\ : Odrv4
    port map (
            O => \N__37400\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7676\ : CascadeMux
    port map (
            O => \N__37391\,
            I => \N__37388\
        );

    \I__7675\ : InMux
    port map (
            O => \N__37388\,
            I => \N__37385\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__37385\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__7673\ : InMux
    port map (
            O => \N__37382\,
            I => \N__37379\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__37379\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__7671\ : InMux
    port map (
            O => \N__37376\,
            I => \N__37373\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__37373\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__7669\ : InMux
    port map (
            O => \N__37370\,
            I => \N__37367\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__37367\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__7667\ : CascadeMux
    port map (
            O => \N__37364\,
            I => \N__37360\
        );

    \I__7666\ : InMux
    port map (
            O => \N__37363\,
            I => \N__37355\
        );

    \I__7665\ : InMux
    port map (
            O => \N__37360\,
            I => \N__37355\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__37355\,
            I => \N__37352\
        );

    \I__7663\ : Odrv4
    port map (
            O => \N__37352\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\
        );

    \I__7662\ : CascadeMux
    port map (
            O => \N__37349\,
            I => \N__37346\
        );

    \I__7661\ : InMux
    port map (
            O => \N__37346\,
            I => \N__37342\
        );

    \I__7660\ : CascadeMux
    port map (
            O => \N__37345\,
            I => \N__37339\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__37342\,
            I => \N__37336\
        );

    \I__7658\ : InMux
    port map (
            O => \N__37339\,
            I => \N__37332\
        );

    \I__7657\ : Span4Mux_v
    port map (
            O => \N__37336\,
            I => \N__37329\
        );

    \I__7656\ : InMux
    port map (
            O => \N__37335\,
            I => \N__37326\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__37332\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7654\ : Odrv4
    port map (
            O => \N__37329\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__37326\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7652\ : InMux
    port map (
            O => \N__37319\,
            I => \N__37315\
        );

    \I__7651\ : InMux
    port map (
            O => \N__37318\,
            I => \N__37312\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__37315\,
            I => \N__37309\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__37312\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__7648\ : Odrv4
    port map (
            O => \N__37309\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__7647\ : InMux
    port map (
            O => \N__37304\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__7646\ : InMux
    port map (
            O => \N__37301\,
            I => \N__37297\
        );

    \I__7645\ : InMux
    port map (
            O => \N__37300\,
            I => \N__37294\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__37297\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__37294\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7642\ : InMux
    port map (
            O => \N__37289\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__7641\ : CascadeMux
    port map (
            O => \N__37286\,
            I => \N__37283\
        );

    \I__7640\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37280\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__37280\,
            I => \N__37277\
        );

    \I__7638\ : Odrv4
    port map (
            O => \N__37277\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__7637\ : CascadeMux
    port map (
            O => \N__37274\,
            I => \N__37271\
        );

    \I__7636\ : InMux
    port map (
            O => \N__37271\,
            I => \N__37268\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__37268\,
            I => \N__37265\
        );

    \I__7634\ : Odrv4
    port map (
            O => \N__37265\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__7633\ : CascadeMux
    port map (
            O => \N__37262\,
            I => \N__37259\
        );

    \I__7632\ : InMux
    port map (
            O => \N__37259\,
            I => \N__37256\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__37256\,
            I => \N__37253\
        );

    \I__7630\ : Odrv4
    port map (
            O => \N__37253\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\
        );

    \I__7629\ : InMux
    port map (
            O => \N__37250\,
            I => \N__37247\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__37247\,
            I => \N__37244\
        );

    \I__7627\ : Odrv4
    port map (
            O => \N__37244\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__7626\ : InMux
    port map (
            O => \N__37241\,
            I => \N__37238\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__37238\,
            I => \N__37235\
        );

    \I__7624\ : Odrv4
    port map (
            O => \N__37235\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__7623\ : InMux
    port map (
            O => \N__37232\,
            I => \N__37229\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__37229\,
            I => \N__37226\
        );

    \I__7621\ : Odrv4
    port map (
            O => \N__37226\,
            I => \current_shift_inst.control_input_axb_19\
        );

    \I__7620\ : InMux
    port map (
            O => \N__37223\,
            I => \N__37220\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__37220\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__7618\ : InMux
    port map (
            O => \N__37217\,
            I => \N__37214\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__37214\,
            I => \N__37211\
        );

    \I__7616\ : Odrv12
    port map (
            O => \N__37211\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\
        );

    \I__7615\ : InMux
    port map (
            O => \N__37208\,
            I => \N__37205\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__37205\,
            I => \N__37202\
        );

    \I__7613\ : Odrv4
    port map (
            O => \N__37202\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__7612\ : InMux
    port map (
            O => \N__37199\,
            I => \N__37196\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__37196\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__7610\ : InMux
    port map (
            O => \N__37193\,
            I => \bfn_14_18_0_\
        );

    \I__7609\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37187\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__37187\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__7607\ : InMux
    port map (
            O => \N__37184\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__7606\ : InMux
    port map (
            O => \N__37181\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__7605\ : InMux
    port map (
            O => \N__37178\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__7604\ : InMux
    port map (
            O => \N__37175\,
            I => \N__37172\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__37172\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__7602\ : InMux
    port map (
            O => \N__37169\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__7601\ : InMux
    port map (
            O => \N__37166\,
            I => \N__37163\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__37163\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__7599\ : InMux
    port map (
            O => \N__37160\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__7598\ : InMux
    port map (
            O => \N__37157\,
            I => \N__37154\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__37154\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__7596\ : InMux
    port map (
            O => \N__37151\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__7595\ : InMux
    port map (
            O => \N__37148\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__7594\ : InMux
    port map (
            O => \N__37145\,
            I => \N__37142\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__37142\,
            I => \N__37139\
        );

    \I__7592\ : Span4Mux_h
    port map (
            O => \N__37139\,
            I => \N__37136\
        );

    \I__7591\ : Odrv4
    port map (
            O => \N__37136\,
            I => \current_shift_inst.control_input_axb_28\
        );

    \I__7590\ : InMux
    port map (
            O => \N__37133\,
            I => \N__37130\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__37130\,
            I => \N__37127\
        );

    \I__7588\ : Odrv12
    port map (
            O => \N__37127\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\
        );

    \I__7587\ : InMux
    port map (
            O => \N__37124\,
            I => \bfn_14_17_0_\
        );

    \I__7586\ : InMux
    port map (
            O => \N__37121\,
            I => \current_shift_inst.un38_control_input_cry_16_s0\
        );

    \I__7585\ : InMux
    port map (
            O => \N__37118\,
            I => \current_shift_inst.un38_control_input_cry_17_s0\
        );

    \I__7584\ : InMux
    port map (
            O => \N__37115\,
            I => \N__37112\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__37112\,
            I => \current_shift_inst.un38_control_input_0_s0_19\
        );

    \I__7582\ : InMux
    port map (
            O => \N__37109\,
            I => \current_shift_inst.un38_control_input_cry_18_s0\
        );

    \I__7581\ : InMux
    port map (
            O => \N__37106\,
            I => \N__37103\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__37103\,
            I => \N__37100\
        );

    \I__7579\ : Odrv4
    port map (
            O => \N__37100\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__7578\ : InMux
    port map (
            O => \N__37097\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__7577\ : InMux
    port map (
            O => \N__37094\,
            I => \N__37091\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__37091\,
            I => \N__37088\
        );

    \I__7575\ : Sp12to4
    port map (
            O => \N__37088\,
            I => \N__37085\
        );

    \I__7574\ : Odrv12
    port map (
            O => \N__37085\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__7573\ : InMux
    port map (
            O => \N__37082\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__7572\ : InMux
    port map (
            O => \N__37079\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__7571\ : InMux
    port map (
            O => \N__37076\,
            I => \N__37073\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__37073\,
            I => \N__37070\
        );

    \I__7569\ : Odrv4
    port map (
            O => \N__37070\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__7568\ : InMux
    port map (
            O => \N__37067\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__7567\ : InMux
    port map (
            O => \N__37064\,
            I => \N__37061\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__37061\,
            I => \N__37058\
        );

    \I__7565\ : Span4Mux_h
    port map (
            O => \N__37058\,
            I => \N__37055\
        );

    \I__7564\ : Odrv4
    port map (
            O => \N__37055\,
            I => \current_shift_inst.un38_control_input_0_s0_7\
        );

    \I__7563\ : InMux
    port map (
            O => \N__37052\,
            I => \current_shift_inst.un38_control_input_cry_6_s0\
        );

    \I__7562\ : InMux
    port map (
            O => \N__37049\,
            I => \N__37046\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__37046\,
            I => \N__37043\
        );

    \I__7560\ : Odrv4
    port map (
            O => \N__37043\,
            I => \current_shift_inst.un38_control_input_0_s0_8\
        );

    \I__7559\ : InMux
    port map (
            O => \N__37040\,
            I => \bfn_14_16_0_\
        );

    \I__7558\ : InMux
    port map (
            O => \N__37037\,
            I => \N__37034\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__37034\,
            I => \N__37031\
        );

    \I__7556\ : Odrv4
    port map (
            O => \N__37031\,
            I => \current_shift_inst.un38_control_input_0_s0_9\
        );

    \I__7555\ : InMux
    port map (
            O => \N__37028\,
            I => \current_shift_inst.un38_control_input_cry_8_s0\
        );

    \I__7554\ : InMux
    port map (
            O => \N__37025\,
            I => \N__37022\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__37022\,
            I => \current_shift_inst.un38_control_input_0_s0_10\
        );

    \I__7552\ : InMux
    port map (
            O => \N__37019\,
            I => \current_shift_inst.un38_control_input_cry_9_s0\
        );

    \I__7551\ : InMux
    port map (
            O => \N__37016\,
            I => \N__37013\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__37013\,
            I => \N__37010\
        );

    \I__7549\ : Span4Mux_v
    port map (
            O => \N__37010\,
            I => \N__37007\
        );

    \I__7548\ : Odrv4
    port map (
            O => \N__37007\,
            I => \current_shift_inst.un38_control_input_0_s0_11\
        );

    \I__7547\ : InMux
    port map (
            O => \N__37004\,
            I => \current_shift_inst.un38_control_input_cry_10_s0\
        );

    \I__7546\ : InMux
    port map (
            O => \N__37001\,
            I => \N__36998\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__36998\,
            I => \N__36995\
        );

    \I__7544\ : Span4Mux_h
    port map (
            O => \N__36995\,
            I => \N__36992\
        );

    \I__7543\ : Odrv4
    port map (
            O => \N__36992\,
            I => \current_shift_inst.un38_control_input_0_s0_12\
        );

    \I__7542\ : InMux
    port map (
            O => \N__36989\,
            I => \current_shift_inst.un38_control_input_cry_11_s0\
        );

    \I__7541\ : InMux
    port map (
            O => \N__36986\,
            I => \N__36983\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__36983\,
            I => \N__36980\
        );

    \I__7539\ : Odrv4
    port map (
            O => \N__36980\,
            I => \current_shift_inst.un38_control_input_0_s0_13\
        );

    \I__7538\ : InMux
    port map (
            O => \N__36977\,
            I => \current_shift_inst.un38_control_input_cry_12_s0\
        );

    \I__7537\ : InMux
    port map (
            O => \N__36974\,
            I => \current_shift_inst.un38_control_input_cry_13_s0\
        );

    \I__7536\ : InMux
    port map (
            O => \N__36971\,
            I => \current_shift_inst.un38_control_input_cry_14_s0\
        );

    \I__7535\ : CascadeMux
    port map (
            O => \N__36968\,
            I => \N__36965\
        );

    \I__7534\ : InMux
    port map (
            O => \N__36965\,
            I => \N__36962\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__36962\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__7532\ : InMux
    port map (
            O => \N__36959\,
            I => \N__36956\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__36956\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\
        );

    \I__7530\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36950\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__36950\,
            I => \N__36947\
        );

    \I__7528\ : Span4Mux_h
    port map (
            O => \N__36947\,
            I => \N__36944\
        );

    \I__7527\ : Odrv4
    port map (
            O => \N__36944\,
            I => \current_shift_inst.un38_control_input_0_s0_3\
        );

    \I__7526\ : InMux
    port map (
            O => \N__36941\,
            I => \current_shift_inst.un38_control_input_cry_2_s0\
        );

    \I__7525\ : InMux
    port map (
            O => \N__36938\,
            I => \N__36935\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__36935\,
            I => \N__36932\
        );

    \I__7523\ : Odrv4
    port map (
            O => \N__36932\,
            I => \current_shift_inst.un38_control_input_0_s0_4\
        );

    \I__7522\ : InMux
    port map (
            O => \N__36929\,
            I => \current_shift_inst.un38_control_input_cry_3_s0\
        );

    \I__7521\ : InMux
    port map (
            O => \N__36926\,
            I => \N__36923\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__36923\,
            I => \N__36920\
        );

    \I__7519\ : Span4Mux_h
    port map (
            O => \N__36920\,
            I => \N__36917\
        );

    \I__7518\ : Odrv4
    port map (
            O => \N__36917\,
            I => \current_shift_inst.un38_control_input_0_s0_5\
        );

    \I__7517\ : InMux
    port map (
            O => \N__36914\,
            I => \current_shift_inst.un38_control_input_cry_4_s0\
        );

    \I__7516\ : InMux
    port map (
            O => \N__36911\,
            I => \N__36908\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__36908\,
            I => \N__36905\
        );

    \I__7514\ : Odrv4
    port map (
            O => \N__36905\,
            I => \current_shift_inst.un38_control_input_0_s0_6\
        );

    \I__7513\ : InMux
    port map (
            O => \N__36902\,
            I => \current_shift_inst.un38_control_input_cry_5_s0\
        );

    \I__7512\ : InMux
    port map (
            O => \N__36899\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__7511\ : InMux
    port map (
            O => \N__36896\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__7510\ : InMux
    port map (
            O => \N__36893\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__7509\ : InMux
    port map (
            O => \N__36890\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__7508\ : InMux
    port map (
            O => \N__36887\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__7507\ : InMux
    port map (
            O => \N__36884\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__7506\ : IoInMux
    port map (
            O => \N__36881\,
            I => \N__36871\
        );

    \I__7505\ : InMux
    port map (
            O => \N__36880\,
            I => \N__36844\
        );

    \I__7504\ : InMux
    port map (
            O => \N__36879\,
            I => \N__36844\
        );

    \I__7503\ : InMux
    port map (
            O => \N__36878\,
            I => \N__36844\
        );

    \I__7502\ : InMux
    port map (
            O => \N__36877\,
            I => \N__36835\
        );

    \I__7501\ : InMux
    port map (
            O => \N__36876\,
            I => \N__36835\
        );

    \I__7500\ : InMux
    port map (
            O => \N__36875\,
            I => \N__36835\
        );

    \I__7499\ : InMux
    port map (
            O => \N__36874\,
            I => \N__36835\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__36871\,
            I => \N__36828\
        );

    \I__7497\ : InMux
    port map (
            O => \N__36870\,
            I => \N__36819\
        );

    \I__7496\ : InMux
    port map (
            O => \N__36869\,
            I => \N__36819\
        );

    \I__7495\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36819\
        );

    \I__7494\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36819\
        );

    \I__7493\ : InMux
    port map (
            O => \N__36866\,
            I => \N__36810\
        );

    \I__7492\ : InMux
    port map (
            O => \N__36865\,
            I => \N__36810\
        );

    \I__7491\ : InMux
    port map (
            O => \N__36864\,
            I => \N__36810\
        );

    \I__7490\ : InMux
    port map (
            O => \N__36863\,
            I => \N__36810\
        );

    \I__7489\ : InMux
    port map (
            O => \N__36862\,
            I => \N__36801\
        );

    \I__7488\ : InMux
    port map (
            O => \N__36861\,
            I => \N__36801\
        );

    \I__7487\ : InMux
    port map (
            O => \N__36860\,
            I => \N__36801\
        );

    \I__7486\ : InMux
    port map (
            O => \N__36859\,
            I => \N__36801\
        );

    \I__7485\ : InMux
    port map (
            O => \N__36858\,
            I => \N__36792\
        );

    \I__7484\ : InMux
    port map (
            O => \N__36857\,
            I => \N__36792\
        );

    \I__7483\ : InMux
    port map (
            O => \N__36856\,
            I => \N__36792\
        );

    \I__7482\ : InMux
    port map (
            O => \N__36855\,
            I => \N__36792\
        );

    \I__7481\ : InMux
    port map (
            O => \N__36854\,
            I => \N__36783\
        );

    \I__7480\ : InMux
    port map (
            O => \N__36853\,
            I => \N__36783\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36852\,
            I => \N__36783\
        );

    \I__7478\ : InMux
    port map (
            O => \N__36851\,
            I => \N__36783\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__36844\,
            I => \N__36778\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__36835\,
            I => \N__36778\
        );

    \I__7475\ : InMux
    port map (
            O => \N__36834\,
            I => \N__36769\
        );

    \I__7474\ : InMux
    port map (
            O => \N__36833\,
            I => \N__36769\
        );

    \I__7473\ : InMux
    port map (
            O => \N__36832\,
            I => \N__36769\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36831\,
            I => \N__36769\
        );

    \I__7471\ : IoSpan4Mux
    port map (
            O => \N__36828\,
            I => \N__36766\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__36819\,
            I => \N__36761\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__36810\,
            I => \N__36761\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__36801\,
            I => \N__36750\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__36792\,
            I => \N__36750\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__36783\,
            I => \N__36750\
        );

    \I__7465\ : Span4Mux_v
    port map (
            O => \N__36778\,
            I => \N__36750\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__36769\,
            I => \N__36750\
        );

    \I__7463\ : Span4Mux_s2_v
    port map (
            O => \N__36766\,
            I => \N__36747\
        );

    \I__7462\ : Span4Mux_v
    port map (
            O => \N__36761\,
            I => \N__36742\
        );

    \I__7461\ : Span4Mux_v
    port map (
            O => \N__36750\,
            I => \N__36742\
        );

    \I__7460\ : Span4Mux_v
    port map (
            O => \N__36747\,
            I => \N__36739\
        );

    \I__7459\ : Span4Mux_h
    port map (
            O => \N__36742\,
            I => \N__36736\
        );

    \I__7458\ : Sp12to4
    port map (
            O => \N__36739\,
            I => \N__36733\
        );

    \I__7457\ : Odrv4
    port map (
            O => \N__36736\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__7456\ : Odrv12
    port map (
            O => \N__36733\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__7455\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36725\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__36725\,
            I => \N__36721\
        );

    \I__7453\ : InMux
    port map (
            O => \N__36724\,
            I => \N__36718\
        );

    \I__7452\ : Span4Mux_h
    port map (
            O => \N__36721\,
            I => \N__36715\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__36718\,
            I => \N__36712\
        );

    \I__7450\ : Span4Mux_h
    port map (
            O => \N__36715\,
            I => \N__36709\
        );

    \I__7449\ : Span12Mux_s10_v
    port map (
            O => \N__36712\,
            I => \N__36706\
        );

    \I__7448\ : Odrv4
    port map (
            O => \N__36709\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__7447\ : Odrv12
    port map (
            O => \N__36706\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__7446\ : CascadeMux
    port map (
            O => \N__36701\,
            I => \N__36697\
        );

    \I__7445\ : InMux
    port map (
            O => \N__36700\,
            I => \N__36693\
        );

    \I__7444\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36689\
        );

    \I__7443\ : InMux
    port map (
            O => \N__36696\,
            I => \N__36686\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__36693\,
            I => \N__36683\
        );

    \I__7441\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36679\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__36689\,
            I => \N__36676\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__36686\,
            I => \N__36673\
        );

    \I__7438\ : Span4Mux_v
    port map (
            O => \N__36683\,
            I => \N__36670\
        );

    \I__7437\ : InMux
    port map (
            O => \N__36682\,
            I => \N__36667\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36679\,
            I => \N__36664\
        );

    \I__7435\ : Span4Mux_h
    port map (
            O => \N__36676\,
            I => \N__36661\
        );

    \I__7434\ : Span4Mux_h
    port map (
            O => \N__36673\,
            I => \N__36658\
        );

    \I__7433\ : Span4Mux_h
    port map (
            O => \N__36670\,
            I => \N__36655\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__36667\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__7431\ : Odrv4
    port map (
            O => \N__36664\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__7430\ : Odrv4
    port map (
            O => \N__36661\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__7429\ : Odrv4
    port map (
            O => \N__36658\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__7428\ : Odrv4
    port map (
            O => \N__36655\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__7427\ : InMux
    port map (
            O => \N__36644\,
            I => \bfn_14_12_0_\
        );

    \I__7426\ : CascadeMux
    port map (
            O => \N__36641\,
            I => \N__36638\
        );

    \I__7425\ : InMux
    port map (
            O => \N__36638\,
            I => \N__36632\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36637\,
            I => \N__36632\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__36632\,
            I => \N__36628\
        );

    \I__7422\ : InMux
    port map (
            O => \N__36631\,
            I => \N__36625\
        );

    \I__7421\ : Span4Mux_h
    port map (
            O => \N__36628\,
            I => \N__36622\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__36625\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7419\ : Odrv4
    port map (
            O => \N__36622\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7418\ : InMux
    port map (
            O => \N__36617\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__7417\ : InMux
    port map (
            O => \N__36614\,
            I => \N__36607\
        );

    \I__7416\ : InMux
    port map (
            O => \N__36613\,
            I => \N__36607\
        );

    \I__7415\ : InMux
    port map (
            O => \N__36612\,
            I => \N__36604\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__36607\,
            I => \N__36601\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__36604\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7412\ : Odrv4
    port map (
            O => \N__36601\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7411\ : InMux
    port map (
            O => \N__36596\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__7410\ : InMux
    port map (
            O => \N__36593\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__7409\ : InMux
    port map (
            O => \N__36590\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__7408\ : InMux
    port map (
            O => \N__36587\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__7407\ : InMux
    port map (
            O => \N__36584\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__7406\ : InMux
    port map (
            O => \N__36581\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__7405\ : InMux
    port map (
            O => \N__36578\,
            I => \bfn_14_13_0_\
        );

    \I__7404\ : InMux
    port map (
            O => \N__36575\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__7403\ : InMux
    port map (
            O => \N__36572\,
            I => \bfn_14_11_0_\
        );

    \I__7402\ : InMux
    port map (
            O => \N__36569\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__7401\ : InMux
    port map (
            O => \N__36566\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__7400\ : InMux
    port map (
            O => \N__36563\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__7399\ : InMux
    port map (
            O => \N__36560\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__7398\ : InMux
    port map (
            O => \N__36557\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__7397\ : InMux
    port map (
            O => \N__36554\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__7396\ : InMux
    port map (
            O => \N__36551\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__7395\ : InMux
    port map (
            O => \N__36548\,
            I => \N__36545\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__36545\,
            I => \N__36542\
        );

    \I__7393\ : Span4Mux_h
    port map (
            O => \N__36542\,
            I => \N__36539\
        );

    \I__7392\ : Span4Mux_v
    port map (
            O => \N__36539\,
            I => \N__36536\
        );

    \I__7391\ : Span4Mux_h
    port map (
            O => \N__36536\,
            I => \N__36533\
        );

    \I__7390\ : Odrv4
    port map (
            O => \N__36533\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\
        );

    \I__7389\ : InMux
    port map (
            O => \N__36530\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__7388\ : CascadeMux
    port map (
            O => \N__36527\,
            I => \N__36524\
        );

    \I__7387\ : InMux
    port map (
            O => \N__36524\,
            I => \N__36521\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__36521\,
            I => \N__36518\
        );

    \I__7385\ : Span4Mux_h
    port map (
            O => \N__36518\,
            I => \N__36515\
        );

    \I__7384\ : Span4Mux_h
    port map (
            O => \N__36515\,
            I => \N__36512\
        );

    \I__7383\ : Sp12to4
    port map (
            O => \N__36512\,
            I => \N__36509\
        );

    \I__7382\ : Odrv12
    port map (
            O => \N__36509\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30\
        );

    \I__7381\ : InMux
    port map (
            O => \N__36506\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__7380\ : InMux
    port map (
            O => \N__36503\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__7379\ : InMux
    port map (
            O => \N__36500\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__7378\ : InMux
    port map (
            O => \N__36497\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__7377\ : InMux
    port map (
            O => \N__36494\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__7376\ : CascadeMux
    port map (
            O => \N__36491\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\
        );

    \I__7375\ : CascadeMux
    port map (
            O => \N__36488\,
            I => \N__36484\
        );

    \I__7374\ : InMux
    port map (
            O => \N__36487\,
            I => \N__36481\
        );

    \I__7373\ : InMux
    port map (
            O => \N__36484\,
            I => \N__36478\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__36481\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__36478\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__7370\ : CascadeMux
    port map (
            O => \N__36473\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15_cascade_\
        );

    \I__7369\ : InMux
    port map (
            O => \N__36470\,
            I => \N__36467\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__36467\,
            I => \N__36464\
        );

    \I__7367\ : Odrv12
    port map (
            O => \N__36464\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__7366\ : InMux
    port map (
            O => \N__36461\,
            I => \N__36456\
        );

    \I__7365\ : InMux
    port map (
            O => \N__36460\,
            I => \N__36453\
        );

    \I__7364\ : InMux
    port map (
            O => \N__36459\,
            I => \N__36450\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__36456\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__36453\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__36450\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__7360\ : InMux
    port map (
            O => \N__36443\,
            I => \N__36437\
        );

    \I__7359\ : InMux
    port map (
            O => \N__36442\,
            I => \N__36437\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__36437\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__7357\ : InMux
    port map (
            O => \N__36434\,
            I => \N__36430\
        );

    \I__7356\ : InMux
    port map (
            O => \N__36433\,
            I => \N__36427\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__36430\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__36427\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__7353\ : CascadeMux
    port map (
            O => \N__36422\,
            I => \N__36419\
        );

    \I__7352\ : InMux
    port map (
            O => \N__36419\,
            I => \N__36413\
        );

    \I__7351\ : InMux
    port map (
            O => \N__36418\,
            I => \N__36413\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__36413\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__7349\ : InMux
    port map (
            O => \N__36410\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30\
        );

    \I__7348\ : CascadeMux
    port map (
            O => \N__36407\,
            I => \N__36404\
        );

    \I__7347\ : InMux
    port map (
            O => \N__36404\,
            I => \N__36401\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__36401\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt26\
        );

    \I__7345\ : InMux
    port map (
            O => \N__36398\,
            I => \N__36392\
        );

    \I__7344\ : InMux
    port map (
            O => \N__36397\,
            I => \N__36392\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__36392\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\
        );

    \I__7342\ : InMux
    port map (
            O => \N__36389\,
            I => \N__36386\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__36386\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\
        );

    \I__7340\ : InMux
    port map (
            O => \N__36383\,
            I => \N__36379\
        );

    \I__7339\ : InMux
    port map (
            O => \N__36382\,
            I => \N__36376\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__36379\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__36376\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\
        );

    \I__7336\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36367\
        );

    \I__7335\ : InMux
    port map (
            O => \N__36370\,
            I => \N__36364\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__36367\,
            I => \N__36359\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__36364\,
            I => \N__36359\
        );

    \I__7332\ : Odrv12
    port map (
            O => \N__36359\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\
        );

    \I__7331\ : InMux
    port map (
            O => \N__36356\,
            I => \N__36353\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__36353\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\
        );

    \I__7329\ : InMux
    port map (
            O => \N__36350\,
            I => \N__36347\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__36347\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\
        );

    \I__7327\ : CascadeMux
    port map (
            O => \N__36344\,
            I => \N__36340\
        );

    \I__7326\ : InMux
    port map (
            O => \N__36343\,
            I => \N__36337\
        );

    \I__7325\ : InMux
    port map (
            O => \N__36340\,
            I => \N__36334\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__36337\,
            I => \N__36331\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__36334\,
            I => \N__36328\
        );

    \I__7322\ : Span4Mux_v
    port map (
            O => \N__36331\,
            I => \N__36325\
        );

    \I__7321\ : Odrv4
    port map (
            O => \N__36328\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__7320\ : Odrv4
    port map (
            O => \N__36325\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__7319\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36317\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__36317\,
            I => \N__36313\
        );

    \I__7317\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36310\
        );

    \I__7316\ : Odrv4
    port map (
            O => \N__36313\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__36310\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__7314\ : CascadeMux
    port map (
            O => \N__36305\,
            I => \N__36302\
        );

    \I__7313\ : InMux
    port map (
            O => \N__36302\,
            I => \N__36299\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__36299\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt24\
        );

    \I__7311\ : InMux
    port map (
            O => \N__36296\,
            I => \N__36293\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__36293\,
            I => \N__36289\
        );

    \I__7309\ : InMux
    port map (
            O => \N__36292\,
            I => \N__36286\
        );

    \I__7308\ : Odrv4
    port map (
            O => \N__36289\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__36286\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__7306\ : CascadeMux
    port map (
            O => \N__36281\,
            I => \N__36278\
        );

    \I__7305\ : InMux
    port map (
            O => \N__36278\,
            I => \N__36275\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__36275\,
            I => \N__36272\
        );

    \I__7303\ : Odrv12
    port map (
            O => \N__36272\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt18\
        );

    \I__7302\ : CascadeMux
    port map (
            O => \N__36269\,
            I => \N__36266\
        );

    \I__7301\ : InMux
    port map (
            O => \N__36266\,
            I => \N__36263\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__36263\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__7299\ : CascadeMux
    port map (
            O => \N__36260\,
            I => \N__36257\
        );

    \I__7298\ : InMux
    port map (
            O => \N__36257\,
            I => \N__36254\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__36254\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt20\
        );

    \I__7296\ : InMux
    port map (
            O => \N__36251\,
            I => \N__36248\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__36248\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\
        );

    \I__7294\ : InMux
    port map (
            O => \N__36245\,
            I => \N__36242\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__36242\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__7292\ : InMux
    port map (
            O => \N__36239\,
            I => \N__36236\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__36236\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__7290\ : CascadeMux
    port map (
            O => \N__36233\,
            I => \N__36230\
        );

    \I__7289\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36227\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__36227\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__7287\ : CascadeMux
    port map (
            O => \N__36224\,
            I => \N__36221\
        );

    \I__7286\ : InMux
    port map (
            O => \N__36221\,
            I => \N__36218\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__36218\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__7284\ : CascadeMux
    port map (
            O => \N__36215\,
            I => \N__36212\
        );

    \I__7283\ : InMux
    port map (
            O => \N__36212\,
            I => \N__36209\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__36209\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__7281\ : CascadeMux
    port map (
            O => \N__36206\,
            I => \N__36203\
        );

    \I__7280\ : InMux
    port map (
            O => \N__36203\,
            I => \N__36200\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__36200\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__7278\ : CascadeMux
    port map (
            O => \N__36197\,
            I => \N__36194\
        );

    \I__7277\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36191\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__36191\,
            I => \N__36188\
        );

    \I__7275\ : Odrv4
    port map (
            O => \N__36188\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__7274\ : CascadeMux
    port map (
            O => \N__36185\,
            I => \N__36182\
        );

    \I__7273\ : InMux
    port map (
            O => \N__36182\,
            I => \N__36179\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__36179\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__7271\ : CascadeMux
    port map (
            O => \N__36176\,
            I => \N__36173\
        );

    \I__7270\ : InMux
    port map (
            O => \N__36173\,
            I => \N__36170\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__36170\,
            I => \N__36167\
        );

    \I__7268\ : Odrv4
    port map (
            O => \N__36167\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__7267\ : CascadeMux
    port map (
            O => \N__36164\,
            I => \N__36161\
        );

    \I__7266\ : InMux
    port map (
            O => \N__36161\,
            I => \N__36158\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__36158\,
            I => \N__36153\
        );

    \I__7264\ : InMux
    port map (
            O => \N__36157\,
            I => \N__36150\
        );

    \I__7263\ : InMux
    port map (
            O => \N__36156\,
            I => \N__36147\
        );

    \I__7262\ : Span4Mux_v
    port map (
            O => \N__36153\,
            I => \N__36140\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__36150\,
            I => \N__36140\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__36147\,
            I => \N__36140\
        );

    \I__7259\ : Span4Mux_v
    port map (
            O => \N__36140\,
            I => \N__36137\
        );

    \I__7258\ : Span4Mux_v
    port map (
            O => \N__36137\,
            I => \N__36134\
        );

    \I__7257\ : Span4Mux_v
    port map (
            O => \N__36134\,
            I => \N__36131\
        );

    \I__7256\ : Odrv4
    port map (
            O => \N__36131\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__7255\ : InMux
    port map (
            O => \N__36128\,
            I => \N__36125\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__36125\,
            I => \N__36121\
        );

    \I__7253\ : InMux
    port map (
            O => \N__36124\,
            I => \N__36118\
        );

    \I__7252\ : Span4Mux_v
    port map (
            O => \N__36121\,
            I => \N__36113\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__36118\,
            I => \N__36113\
        );

    \I__7250\ : Span4Mux_v
    port map (
            O => \N__36113\,
            I => \N__36110\
        );

    \I__7249\ : Span4Mux_v
    port map (
            O => \N__36110\,
            I => \N__36105\
        );

    \I__7248\ : InMux
    port map (
            O => \N__36109\,
            I => \N__36100\
        );

    \I__7247\ : InMux
    port map (
            O => \N__36108\,
            I => \N__36100\
        );

    \I__7246\ : Span4Mux_v
    port map (
            O => \N__36105\,
            I => \N__36097\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__36100\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__7244\ : Odrv4
    port map (
            O => \N__36097\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__7243\ : ClkMux
    port map (
            O => \N__36092\,
            I => \N__36089\
        );

    \I__7242\ : GlobalMux
    port map (
            O => \N__36089\,
            I => \N__36086\
        );

    \I__7241\ : gio2CtrlBuf
    port map (
            O => \N__36086\,
            I => delay_hc_input_c_g
        );

    \I__7240\ : CascadeMux
    port map (
            O => \N__36083\,
            I => \N__36080\
        );

    \I__7239\ : InMux
    port map (
            O => \N__36080\,
            I => \N__36077\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__36077\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__7237\ : CascadeMux
    port map (
            O => \N__36074\,
            I => \N__36071\
        );

    \I__7236\ : InMux
    port map (
            O => \N__36071\,
            I => \N__36068\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__36068\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__7234\ : InMux
    port map (
            O => \N__36065\,
            I => \N__36062\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__36062\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__7232\ : CascadeMux
    port map (
            O => \N__36059\,
            I => \N__36056\
        );

    \I__7231\ : InMux
    port map (
            O => \N__36056\,
            I => \N__36053\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__36053\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__7229\ : CascadeMux
    port map (
            O => \N__36050\,
            I => \N__36047\
        );

    \I__7228\ : InMux
    port map (
            O => \N__36047\,
            I => \N__36044\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__36044\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__7226\ : InMux
    port map (
            O => \N__36041\,
            I => \N__36038\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__36038\,
            I => \N__36035\
        );

    \I__7224\ : Odrv4
    port map (
            O => \N__36035\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__7223\ : CascadeMux
    port map (
            O => \N__36032\,
            I => \N__36029\
        );

    \I__7222\ : InMux
    port map (
            O => \N__36029\,
            I => \N__36026\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__36026\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__7220\ : CascadeMux
    port map (
            O => \N__36023\,
            I => \N__36020\
        );

    \I__7219\ : InMux
    port map (
            O => \N__36020\,
            I => \N__36017\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__36017\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__7217\ : InMux
    port map (
            O => \N__36014\,
            I => \N__36011\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__36011\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__7215\ : InMux
    port map (
            O => \N__36008\,
            I => \N__36005\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__36005\,
            I => \current_shift_inst.control_input_axb_25\
        );

    \I__7213\ : InMux
    port map (
            O => \N__36002\,
            I => \N__35999\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__35999\,
            I => \current_shift_inst.control_input_axb_29\
        );

    \I__7211\ : InMux
    port map (
            O => \N__35996\,
            I => \N__35991\
        );

    \I__7210\ : InMux
    port map (
            O => \N__35995\,
            I => \N__35988\
        );

    \I__7209\ : InMux
    port map (
            O => \N__35994\,
            I => \N__35985\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__35991\,
            I => \N__35982\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__35988\,
            I => \N__35977\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__35985\,
            I => \N__35977\
        );

    \I__7205\ : Span4Mux_h
    port map (
            O => \N__35982\,
            I => \N__35974\
        );

    \I__7204\ : Span4Mux_h
    port map (
            O => \N__35977\,
            I => \N__35971\
        );

    \I__7203\ : Odrv4
    port map (
            O => \N__35974\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7202\ : Odrv4
    port map (
            O => \N__35971\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7201\ : InMux
    port map (
            O => \N__35966\,
            I => \N__35962\
        );

    \I__7200\ : InMux
    port map (
            O => \N__35965\,
            I => \N__35959\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__35962\,
            I => \N__35954\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__35959\,
            I => \N__35951\
        );

    \I__7197\ : InMux
    port map (
            O => \N__35958\,
            I => \N__35946\
        );

    \I__7196\ : InMux
    port map (
            O => \N__35957\,
            I => \N__35946\
        );

    \I__7195\ : Span4Mux_v
    port map (
            O => \N__35954\,
            I => \N__35943\
        );

    \I__7194\ : Span4Mux_h
    port map (
            O => \N__35951\,
            I => \N__35940\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__35946\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7192\ : Odrv4
    port map (
            O => \N__35943\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7191\ : Odrv4
    port map (
            O => \N__35940\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7190\ : ClkMux
    port map (
            O => \N__35933\,
            I => \N__35930\
        );

    \I__7189\ : GlobalMux
    port map (
            O => \N__35930\,
            I => \N__35927\
        );

    \I__7188\ : gio2CtrlBuf
    port map (
            O => \N__35927\,
            I => delay_tr_input_c_g
        );

    \I__7187\ : IoInMux
    port map (
            O => \N__35924\,
            I => \N__35921\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__35921\,
            I => \N__35918\
        );

    \I__7185\ : Span4Mux_s0_v
    port map (
            O => \N__35918\,
            I => \N__35915\
        );

    \I__7184\ : Span4Mux_v
    port map (
            O => \N__35915\,
            I => \N__35912\
        );

    \I__7183\ : Span4Mux_v
    port map (
            O => \N__35912\,
            I => \N__35907\
        );

    \I__7182\ : InMux
    port map (
            O => \N__35911\,
            I => \N__35904\
        );

    \I__7181\ : InMux
    port map (
            O => \N__35910\,
            I => \N__35901\
        );

    \I__7180\ : Odrv4
    port map (
            O => \N__35907\,
            I => s1_phy_c
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__35904\,
            I => s1_phy_c
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__35901\,
            I => s1_phy_c
        );

    \I__7177\ : InMux
    port map (
            O => \N__35894\,
            I => \N__35891\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__35891\,
            I => \N__35883\
        );

    \I__7175\ : InMux
    port map (
            O => \N__35890\,
            I => \N__35878\
        );

    \I__7174\ : InMux
    port map (
            O => \N__35889\,
            I => \N__35878\
        );

    \I__7173\ : InMux
    port map (
            O => \N__35888\,
            I => \N__35875\
        );

    \I__7172\ : CascadeMux
    port map (
            O => \N__35887\,
            I => \N__35871\
        );

    \I__7171\ : InMux
    port map (
            O => \N__35886\,
            I => \N__35868\
        );

    \I__7170\ : Span4Mux_v
    port map (
            O => \N__35883\,
            I => \N__35863\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__35878\,
            I => \N__35863\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__35875\,
            I => \N__35860\
        );

    \I__7167\ : InMux
    port map (
            O => \N__35874\,
            I => \N__35857\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35871\,
            I => \N__35854\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__35868\,
            I => \N__35851\
        );

    \I__7164\ : Span4Mux_v
    port map (
            O => \N__35863\,
            I => \N__35848\
        );

    \I__7163\ : Span4Mux_v
    port map (
            O => \N__35860\,
            I => \N__35845\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__35857\,
            I => state_3
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__35854\,
            I => state_3
        );

    \I__7160\ : Odrv12
    port map (
            O => \N__35851\,
            I => state_3
        );

    \I__7159\ : Odrv4
    port map (
            O => \N__35848\,
            I => state_3
        );

    \I__7158\ : Odrv4
    port map (
            O => \N__35845\,
            I => state_3
        );

    \I__7157\ : IoInMux
    port map (
            O => \N__35834\,
            I => \N__35831\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__35831\,
            I => \N__35828\
        );

    \I__7155\ : Odrv12
    port map (
            O => \N__35828\,
            I => \current_shift_inst.timer_s1.N_161_i\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35825\,
            I => \N__35821\
        );

    \I__7153\ : InMux
    port map (
            O => \N__35824\,
            I => \N__35818\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__35821\,
            I => \N__35815\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__35818\,
            I => \N__35811\
        );

    \I__7150\ : Span4Mux_v
    port map (
            O => \N__35815\,
            I => \N__35808\
        );

    \I__7149\ : InMux
    port map (
            O => \N__35814\,
            I => \N__35805\
        );

    \I__7148\ : Span12Mux_s6_v
    port map (
            O => \N__35811\,
            I => \N__35802\
        );

    \I__7147\ : Span4Mux_v
    port map (
            O => \N__35808\,
            I => \N__35799\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__35805\,
            I => \N__35795\
        );

    \I__7145\ : Span12Mux_v
    port map (
            O => \N__35802\,
            I => \N__35792\
        );

    \I__7144\ : Span4Mux_v
    port map (
            O => \N__35799\,
            I => \N__35789\
        );

    \I__7143\ : InMux
    port map (
            O => \N__35798\,
            I => \N__35786\
        );

    \I__7142\ : Span4Mux_h
    port map (
            O => \N__35795\,
            I => \N__35783\
        );

    \I__7141\ : Odrv12
    port map (
            O => \N__35792\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7140\ : Odrv4
    port map (
            O => \N__35789\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__35786\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7138\ : Odrv4
    port map (
            O => \N__35783\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7137\ : IoInMux
    port map (
            O => \N__35774\,
            I => \N__35771\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__35771\,
            I => \N__35768\
        );

    \I__7135\ : Odrv4
    port map (
            O => \N__35768\,
            I => s2_phy_c
        );

    \I__7134\ : InMux
    port map (
            O => \N__35765\,
            I => \N__35762\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__35762\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__7132\ : InMux
    port map (
            O => \N__35759\,
            I => \N__35756\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__35756\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__7130\ : InMux
    port map (
            O => \N__35753\,
            I => \N__35750\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__35750\,
            I => \current_shift_inst.control_input_axb_18\
        );

    \I__7128\ : InMux
    port map (
            O => \N__35747\,
            I => \N__35744\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__35744\,
            I => \current_shift_inst.control_input_axb_17\
        );

    \I__7126\ : InMux
    port map (
            O => \N__35741\,
            I => \N__35738\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__35738\,
            I => \current_shift_inst.control_input_axb_20\
        );

    \I__7124\ : InMux
    port map (
            O => \N__35735\,
            I => \N__35732\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__35732\,
            I => \current_shift_inst.control_input_axb_21\
        );

    \I__7122\ : InMux
    port map (
            O => \N__35729\,
            I => \N__35726\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__35726\,
            I => \current_shift_inst.control_input_axb_22\
        );

    \I__7120\ : InMux
    port map (
            O => \N__35723\,
            I => \N__35720\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__35720\,
            I => \current_shift_inst.control_input_axb_27\
        );

    \I__7118\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35714\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__35714\,
            I => \current_shift_inst.control_input_axb_26\
        );

    \I__7116\ : InMux
    port map (
            O => \N__35711\,
            I => \N__35708\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__35708\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__7114\ : InMux
    port map (
            O => \N__35705\,
            I => \N__35701\
        );

    \I__7113\ : InMux
    port map (
            O => \N__35704\,
            I => \N__35696\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__35701\,
            I => \N__35693\
        );

    \I__7111\ : InMux
    port map (
            O => \N__35700\,
            I => \N__35690\
        );

    \I__7110\ : InMux
    port map (
            O => \N__35699\,
            I => \N__35687\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__35696\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__7108\ : Odrv4
    port map (
            O => \N__35693\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__35690\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__35687\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35678\,
            I => \N__35675\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__35675\,
            I => \N__35672\
        );

    \I__7103\ : Span4Mux_v
    port map (
            O => \N__35672\,
            I => \N__35668\
        );

    \I__7102\ : InMux
    port map (
            O => \N__35671\,
            I => \N__35664\
        );

    \I__7101\ : Span4Mux_v
    port map (
            O => \N__35668\,
            I => \N__35660\
        );

    \I__7100\ : InMux
    port map (
            O => \N__35667\,
            I => \N__35657\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__35664\,
            I => \N__35654\
        );

    \I__7098\ : InMux
    port map (
            O => \N__35663\,
            I => \N__35651\
        );

    \I__7097\ : Span4Mux_v
    port map (
            O => \N__35660\,
            I => \N__35646\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__35657\,
            I => \N__35646\
        );

    \I__7095\ : Span12Mux_h
    port map (
            O => \N__35654\,
            I => \N__35643\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__35651\,
            I => \N__35640\
        );

    \I__7093\ : Span4Mux_v
    port map (
            O => \N__35646\,
            I => \N__35637\
        );

    \I__7092\ : Span12Mux_v
    port map (
            O => \N__35643\,
            I => \N__35634\
        );

    \I__7091\ : Span12Mux_h
    port map (
            O => \N__35640\,
            I => \N__35631\
        );

    \I__7090\ : Span4Mux_h
    port map (
            O => \N__35637\,
            I => \N__35628\
        );

    \I__7089\ : Odrv12
    port map (
            O => \N__35634\,
            I => il_max_comp1_c
        );

    \I__7088\ : Odrv12
    port map (
            O => \N__35631\,
            I => il_max_comp1_c
        );

    \I__7087\ : Odrv4
    port map (
            O => \N__35628\,
            I => il_max_comp1_c
        );

    \I__7086\ : IoInMux
    port map (
            O => \N__35621\,
            I => \N__35618\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__35618\,
            I => \N__35615\
        );

    \I__7084\ : Span4Mux_s1_v
    port map (
            O => \N__35615\,
            I => \N__35612\
        );

    \I__7083\ : Sp12to4
    port map (
            O => \N__35612\,
            I => \N__35609\
        );

    \I__7082\ : Span12Mux_h
    port map (
            O => \N__35609\,
            I => \N__35606\
        );

    \I__7081\ : Span12Mux_v
    port map (
            O => \N__35606\,
            I => \N__35602\
        );

    \I__7080\ : InMux
    port map (
            O => \N__35605\,
            I => \N__35599\
        );

    \I__7079\ : Odrv12
    port map (
            O => \N__35602\,
            I => test_c
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__35599\,
            I => test_c
        );

    \I__7077\ : InMux
    port map (
            O => \N__35594\,
            I => \N__35591\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__35591\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__7075\ : InMux
    port map (
            O => \N__35588\,
            I => \N__35585\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__35585\,
            I => \current_shift_inst.control_input_axb_16\
        );

    \I__7073\ : InMux
    port map (
            O => \N__35582\,
            I => \N__35579\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__35579\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__7071\ : InMux
    port map (
            O => \N__35576\,
            I => \N__35573\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__35573\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__7069\ : InMux
    port map (
            O => \N__35570\,
            I => \N__35567\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__35567\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__7067\ : InMux
    port map (
            O => \N__35564\,
            I => \N__35561\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__35561\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__7065\ : CascadeMux
    port map (
            O => \N__35558\,
            I => \N__35554\
        );

    \I__7064\ : CascadeMux
    port map (
            O => \N__35557\,
            I => \N__35551\
        );

    \I__7063\ : InMux
    port map (
            O => \N__35554\,
            I => \N__35546\
        );

    \I__7062\ : InMux
    port map (
            O => \N__35551\,
            I => \N__35546\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__35546\,
            I => \N__35542\
        );

    \I__7060\ : InMux
    port map (
            O => \N__35545\,
            I => \N__35539\
        );

    \I__7059\ : Span4Mux_h
    port map (
            O => \N__35542\,
            I => \N__35536\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__35539\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__7057\ : Odrv4
    port map (
            O => \N__35536\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__7056\ : InMux
    port map (
            O => \N__35531\,
            I => \N__35528\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__35528\,
            I => \N__35522\
        );

    \I__7054\ : InMux
    port map (
            O => \N__35527\,
            I => \N__35519\
        );

    \I__7053\ : CascadeMux
    port map (
            O => \N__35526\,
            I => \N__35516\
        );

    \I__7052\ : InMux
    port map (
            O => \N__35525\,
            I => \N__35513\
        );

    \I__7051\ : Span4Mux_v
    port map (
            O => \N__35522\,
            I => \N__35508\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__35519\,
            I => \N__35508\
        );

    \I__7049\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35505\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__35513\,
            I => \N__35502\
        );

    \I__7047\ : Span4Mux_h
    port map (
            O => \N__35508\,
            I => \N__35499\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__35505\,
            I => \N__35496\
        );

    \I__7045\ : Span4Mux_v
    port map (
            O => \N__35502\,
            I => \N__35493\
        );

    \I__7044\ : Span4Mux_v
    port map (
            O => \N__35499\,
            I => \N__35488\
        );

    \I__7043\ : Span4Mux_v
    port map (
            O => \N__35496\,
            I => \N__35488\
        );

    \I__7042\ : Odrv4
    port map (
            O => \N__35493\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__7041\ : Odrv4
    port map (
            O => \N__35488\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__7040\ : InMux
    port map (
            O => \N__35483\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__7039\ : CascadeMux
    port map (
            O => \N__35480\,
            I => \N__35476\
        );

    \I__7038\ : CascadeMux
    port map (
            O => \N__35479\,
            I => \N__35473\
        );

    \I__7037\ : InMux
    port map (
            O => \N__35476\,
            I => \N__35470\
        );

    \I__7036\ : InMux
    port map (
            O => \N__35473\,
            I => \N__35467\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__35470\,
            I => \N__35464\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__35467\,
            I => \N__35460\
        );

    \I__7033\ : Span4Mux_h
    port map (
            O => \N__35464\,
            I => \N__35457\
        );

    \I__7032\ : InMux
    port map (
            O => \N__35463\,
            I => \N__35454\
        );

    \I__7031\ : Span4Mux_v
    port map (
            O => \N__35460\,
            I => \N__35451\
        );

    \I__7030\ : Span4Mux_h
    port map (
            O => \N__35457\,
            I => \N__35448\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__35454\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__7028\ : Odrv4
    port map (
            O => \N__35451\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__7027\ : Odrv4
    port map (
            O => \N__35448\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__7026\ : InMux
    port map (
            O => \N__35441\,
            I => \N__35437\
        );

    \I__7025\ : InMux
    port map (
            O => \N__35440\,
            I => \N__35434\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__35437\,
            I => \N__35431\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__35434\,
            I => \N__35426\
        );

    \I__7022\ : Span4Mux_v
    port map (
            O => \N__35431\,
            I => \N__35423\
        );

    \I__7021\ : InMux
    port map (
            O => \N__35430\,
            I => \N__35418\
        );

    \I__7020\ : InMux
    port map (
            O => \N__35429\,
            I => \N__35418\
        );

    \I__7019\ : Span4Mux_v
    port map (
            O => \N__35426\,
            I => \N__35415\
        );

    \I__7018\ : Sp12to4
    port map (
            O => \N__35423\,
            I => \N__35410\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__35418\,
            I => \N__35410\
        );

    \I__7016\ : Span4Mux_v
    port map (
            O => \N__35415\,
            I => \N__35407\
        );

    \I__7015\ : Odrv12
    port map (
            O => \N__35410\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__7014\ : Odrv4
    port map (
            O => \N__35407\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__7013\ : InMux
    port map (
            O => \N__35402\,
            I => \bfn_13_13_0_\
        );

    \I__7012\ : InMux
    port map (
            O => \N__35399\,
            I => \N__35395\
        );

    \I__7011\ : InMux
    port map (
            O => \N__35398\,
            I => \N__35392\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__35395\,
            I => \N__35386\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__35392\,
            I => \N__35386\
        );

    \I__7008\ : InMux
    port map (
            O => \N__35391\,
            I => \N__35383\
        );

    \I__7007\ : Span4Mux_v
    port map (
            O => \N__35386\,
            I => \N__35380\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__35383\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__7005\ : Odrv4
    port map (
            O => \N__35380\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__7004\ : InMux
    port map (
            O => \N__35375\,
            I => \N__35371\
        );

    \I__7003\ : InMux
    port map (
            O => \N__35374\,
            I => \N__35367\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__35371\,
            I => \N__35364\
        );

    \I__7001\ : InMux
    port map (
            O => \N__35370\,
            I => \N__35360\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__35367\,
            I => \N__35357\
        );

    \I__6999\ : Span4Mux_v
    port map (
            O => \N__35364\,
            I => \N__35354\
        );

    \I__6998\ : InMux
    port map (
            O => \N__35363\,
            I => \N__35351\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__35360\,
            I => \N__35348\
        );

    \I__6996\ : Span4Mux_v
    port map (
            O => \N__35357\,
            I => \N__35345\
        );

    \I__6995\ : Span4Mux_v
    port map (
            O => \N__35354\,
            I => \N__35342\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__35351\,
            I => \N__35337\
        );

    \I__6993\ : Span12Mux_v
    port map (
            O => \N__35348\,
            I => \N__35337\
        );

    \I__6992\ : Span4Mux_h
    port map (
            O => \N__35345\,
            I => \N__35334\
        );

    \I__6991\ : Span4Mux_h
    port map (
            O => \N__35342\,
            I => \N__35331\
        );

    \I__6990\ : Odrv12
    port map (
            O => \N__35337\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__6989\ : Odrv4
    port map (
            O => \N__35334\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__6988\ : Odrv4
    port map (
            O => \N__35331\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__6987\ : InMux
    port map (
            O => \N__35324\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__6986\ : InMux
    port map (
            O => \N__35321\,
            I => \N__35318\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__35318\,
            I => \N__35314\
        );

    \I__6984\ : InMux
    port map (
            O => \N__35317\,
            I => \N__35311\
        );

    \I__6983\ : Span4Mux_h
    port map (
            O => \N__35314\,
            I => \N__35308\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__35311\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__6981\ : Odrv4
    port map (
            O => \N__35308\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__6980\ : CascadeMux
    port map (
            O => \N__35303\,
            I => \N__35300\
        );

    \I__6979\ : InMux
    port map (
            O => \N__35300\,
            I => \N__35296\
        );

    \I__6978\ : InMux
    port map (
            O => \N__35299\,
            I => \N__35293\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__35296\,
            I => \N__35287\
        );

    \I__6976\ : LocalMux
    port map (
            O => \N__35293\,
            I => \N__35287\
        );

    \I__6975\ : InMux
    port map (
            O => \N__35292\,
            I => \N__35284\
        );

    \I__6974\ : Span4Mux_h
    port map (
            O => \N__35287\,
            I => \N__35281\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__35284\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__6972\ : Odrv4
    port map (
            O => \N__35281\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__6971\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35272\
        );

    \I__6970\ : InMux
    port map (
            O => \N__35275\,
            I => \N__35267\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__35272\,
            I => \N__35264\
        );

    \I__6968\ : InMux
    port map (
            O => \N__35271\,
            I => \N__35259\
        );

    \I__6967\ : InMux
    port map (
            O => \N__35270\,
            I => \N__35259\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__35267\,
            I => \N__35256\
        );

    \I__6965\ : Span4Mux_v
    port map (
            O => \N__35264\,
            I => \N__35251\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__35259\,
            I => \N__35251\
        );

    \I__6963\ : Span4Mux_h
    port map (
            O => \N__35256\,
            I => \N__35248\
        );

    \I__6962\ : Span4Mux_h
    port map (
            O => \N__35251\,
            I => \N__35243\
        );

    \I__6961\ : Span4Mux_v
    port map (
            O => \N__35248\,
            I => \N__35243\
        );

    \I__6960\ : Odrv4
    port map (
            O => \N__35243\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__6959\ : InMux
    port map (
            O => \N__35240\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__6958\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35234\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__35234\,
            I => \N__35230\
        );

    \I__6956\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35227\
        );

    \I__6955\ : Span4Mux_h
    port map (
            O => \N__35230\,
            I => \N__35224\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__35227\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__6953\ : Odrv4
    port map (
            O => \N__35224\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__6952\ : CascadeMux
    port map (
            O => \N__35219\,
            I => \N__35215\
        );

    \I__6951\ : CascadeMux
    port map (
            O => \N__35218\,
            I => \N__35212\
        );

    \I__6950\ : InMux
    port map (
            O => \N__35215\,
            I => \N__35207\
        );

    \I__6949\ : InMux
    port map (
            O => \N__35212\,
            I => \N__35207\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__35207\,
            I => \N__35203\
        );

    \I__6947\ : InMux
    port map (
            O => \N__35206\,
            I => \N__35200\
        );

    \I__6946\ : Span4Mux_h
    port map (
            O => \N__35203\,
            I => \N__35197\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__35200\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__6944\ : Odrv4
    port map (
            O => \N__35197\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__6943\ : InMux
    port map (
            O => \N__35192\,
            I => \N__35186\
        );

    \I__6942\ : InMux
    port map (
            O => \N__35191\,
            I => \N__35183\
        );

    \I__6941\ : InMux
    port map (
            O => \N__35190\,
            I => \N__35180\
        );

    \I__6940\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35177\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__35186\,
            I => \N__35170\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__35183\,
            I => \N__35170\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__35180\,
            I => \N__35170\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__35177\,
            I => \N__35167\
        );

    \I__6935\ : Span4Mux_v
    port map (
            O => \N__35170\,
            I => \N__35164\
        );

    \I__6934\ : Span4Mux_h
    port map (
            O => \N__35167\,
            I => \N__35161\
        );

    \I__6933\ : Odrv4
    port map (
            O => \N__35164\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__6932\ : Odrv4
    port map (
            O => \N__35161\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__6931\ : InMux
    port map (
            O => \N__35156\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__6930\ : InMux
    port map (
            O => \N__35153\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__6929\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35144\
        );

    \I__6928\ : InMux
    port map (
            O => \N__35149\,
            I => \N__35141\
        );

    \I__6927\ : InMux
    port map (
            O => \N__35148\,
            I => \N__35138\
        );

    \I__6926\ : InMux
    port map (
            O => \N__35147\,
            I => \N__35135\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__35144\,
            I => \N__35132\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__35141\,
            I => \N__35127\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__35138\,
            I => \N__35127\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__35135\,
            I => \N__35124\
        );

    \I__6921\ : Span4Mux_h
    port map (
            O => \N__35132\,
            I => \N__35121\
        );

    \I__6920\ : Span4Mux_v
    port map (
            O => \N__35127\,
            I => \N__35118\
        );

    \I__6919\ : Span4Mux_h
    port map (
            O => \N__35124\,
            I => \N__35115\
        );

    \I__6918\ : Span4Mux_v
    port map (
            O => \N__35121\,
            I => \N__35112\
        );

    \I__6917\ : Odrv4
    port map (
            O => \N__35118\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__6916\ : Odrv4
    port map (
            O => \N__35115\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__35112\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__6914\ : CEMux
    port map (
            O => \N__35105\,
            I => \N__35101\
        );

    \I__6913\ : CEMux
    port map (
            O => \N__35104\,
            I => \N__35096\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__35101\,
            I => \N__35093\
        );

    \I__6911\ : CEMux
    port map (
            O => \N__35100\,
            I => \N__35090\
        );

    \I__6910\ : CEMux
    port map (
            O => \N__35099\,
            I => \N__35087\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__35096\,
            I => \N__35083\
        );

    \I__6908\ : Span4Mux_v
    port map (
            O => \N__35093\,
            I => \N__35080\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__35090\,
            I => \N__35077\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__35087\,
            I => \N__35074\
        );

    \I__6905\ : CEMux
    port map (
            O => \N__35086\,
            I => \N__35071\
        );

    \I__6904\ : Span4Mux_h
    port map (
            O => \N__35083\,
            I => \N__35068\
        );

    \I__6903\ : Span4Mux_h
    port map (
            O => \N__35080\,
            I => \N__35065\
        );

    \I__6902\ : Span4Mux_h
    port map (
            O => \N__35077\,
            I => \N__35062\
        );

    \I__6901\ : Span4Mux_v
    port map (
            O => \N__35074\,
            I => \N__35059\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__35071\,
            I => \N__35056\
        );

    \I__6899\ : Span4Mux_v
    port map (
            O => \N__35068\,
            I => \N__35053\
        );

    \I__6898\ : Span4Mux_v
    port map (
            O => \N__35065\,
            I => \N__35048\
        );

    \I__6897\ : Span4Mux_v
    port map (
            O => \N__35062\,
            I => \N__35048\
        );

    \I__6896\ : Span4Mux_v
    port map (
            O => \N__35059\,
            I => \N__35043\
        );

    \I__6895\ : Span4Mux_h
    port map (
            O => \N__35056\,
            I => \N__35043\
        );

    \I__6894\ : Odrv4
    port map (
            O => \N__35053\,
            I => \delay_measurement_inst.delay_tr_timer.N_165_i\
        );

    \I__6893\ : Odrv4
    port map (
            O => \N__35048\,
            I => \delay_measurement_inst.delay_tr_timer.N_165_i\
        );

    \I__6892\ : Odrv4
    port map (
            O => \N__35043\,
            I => \delay_measurement_inst.delay_tr_timer.N_165_i\
        );

    \I__6891\ : InMux
    port map (
            O => \N__35036\,
            I => \N__35030\
        );

    \I__6890\ : InMux
    port map (
            O => \N__35035\,
            I => \N__35030\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__35030\,
            I => \N__35026\
        );

    \I__6888\ : InMux
    port map (
            O => \N__35029\,
            I => \N__35023\
        );

    \I__6887\ : Span4Mux_h
    port map (
            O => \N__35026\,
            I => \N__35020\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__35023\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__6885\ : Odrv4
    port map (
            O => \N__35020\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__6884\ : InMux
    port map (
            O => \N__35015\,
            I => \N__35011\
        );

    \I__6883\ : InMux
    port map (
            O => \N__35014\,
            I => \N__35008\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__35011\,
            I => \N__35002\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__35008\,
            I => \N__35002\
        );

    \I__6880\ : InMux
    port map (
            O => \N__35007\,
            I => \N__34999\
        );

    \I__6879\ : Span4Mux_v
    port map (
            O => \N__35002\,
            I => \N__34993\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__34999\,
            I => \N__34993\
        );

    \I__6877\ : InMux
    port map (
            O => \N__34998\,
            I => \N__34990\
        );

    \I__6876\ : Span4Mux_h
    port map (
            O => \N__34993\,
            I => \N__34985\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__34990\,
            I => \N__34985\
        );

    \I__6874\ : Odrv4
    port map (
            O => \N__34985\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__6873\ : InMux
    port map (
            O => \N__34982\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__6872\ : CascadeMux
    port map (
            O => \N__34979\,
            I => \N__34976\
        );

    \I__6871\ : InMux
    port map (
            O => \N__34976\,
            I => \N__34973\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__34973\,
            I => \N__34969\
        );

    \I__6869\ : InMux
    port map (
            O => \N__34972\,
            I => \N__34966\
        );

    \I__6868\ : Span4Mux_v
    port map (
            O => \N__34969\,
            I => \N__34962\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__34966\,
            I => \N__34959\
        );

    \I__6866\ : InMux
    port map (
            O => \N__34965\,
            I => \N__34956\
        );

    \I__6865\ : Span4Mux_h
    port map (
            O => \N__34962\,
            I => \N__34953\
        );

    \I__6864\ : Span4Mux_h
    port map (
            O => \N__34959\,
            I => \N__34950\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__34956\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__6862\ : Odrv4
    port map (
            O => \N__34953\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__6861\ : Odrv4
    port map (
            O => \N__34950\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__6860\ : InMux
    port map (
            O => \N__34943\,
            I => \N__34939\
        );

    \I__6859\ : InMux
    port map (
            O => \N__34942\,
            I => \N__34936\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__34939\,
            I => \N__34931\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__34936\,
            I => \N__34928\
        );

    \I__6856\ : InMux
    port map (
            O => \N__34935\,
            I => \N__34925\
        );

    \I__6855\ : CascadeMux
    port map (
            O => \N__34934\,
            I => \N__34922\
        );

    \I__6854\ : Span4Mux_h
    port map (
            O => \N__34931\,
            I => \N__34919\
        );

    \I__6853\ : Span4Mux_v
    port map (
            O => \N__34928\,
            I => \N__34916\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__34925\,
            I => \N__34913\
        );

    \I__6851\ : InMux
    port map (
            O => \N__34922\,
            I => \N__34910\
        );

    \I__6850\ : Span4Mux_v
    port map (
            O => \N__34919\,
            I => \N__34907\
        );

    \I__6849\ : Span4Mux_h
    port map (
            O => \N__34916\,
            I => \N__34900\
        );

    \I__6848\ : Span4Mux_v
    port map (
            O => \N__34913\,
            I => \N__34900\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__34910\,
            I => \N__34900\
        );

    \I__6846\ : Odrv4
    port map (
            O => \N__34907\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__6845\ : Odrv4
    port map (
            O => \N__34900\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__6844\ : InMux
    port map (
            O => \N__34895\,
            I => \bfn_13_12_0_\
        );

    \I__6843\ : CascadeMux
    port map (
            O => \N__34892\,
            I => \N__34888\
        );

    \I__6842\ : CascadeMux
    port map (
            O => \N__34891\,
            I => \N__34885\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34888\,
            I => \N__34882\
        );

    \I__6840\ : InMux
    port map (
            O => \N__34885\,
            I => \N__34879\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__34882\,
            I => \N__34875\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__34879\,
            I => \N__34872\
        );

    \I__6837\ : InMux
    port map (
            O => \N__34878\,
            I => \N__34869\
        );

    \I__6836\ : Span4Mux_v
    port map (
            O => \N__34875\,
            I => \N__34866\
        );

    \I__6835\ : Span4Mux_h
    port map (
            O => \N__34872\,
            I => \N__34863\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__34869\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__6833\ : Odrv4
    port map (
            O => \N__34866\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__6832\ : Odrv4
    port map (
            O => \N__34863\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__6831\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34853\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__34853\,
            I => \N__34849\
        );

    \I__6829\ : InMux
    port map (
            O => \N__34852\,
            I => \N__34846\
        );

    \I__6828\ : Span4Mux_v
    port map (
            O => \N__34849\,
            I => \N__34840\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__34846\,
            I => \N__34840\
        );

    \I__6826\ : InMux
    port map (
            O => \N__34845\,
            I => \N__34837\
        );

    \I__6825\ : Span4Mux_v
    port map (
            O => \N__34840\,
            I => \N__34834\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__34837\,
            I => \N__34831\
        );

    \I__6823\ : Span4Mux_h
    port map (
            O => \N__34834\,
            I => \N__34825\
        );

    \I__6822\ : Span4Mux_h
    port map (
            O => \N__34831\,
            I => \N__34825\
        );

    \I__6821\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34822\
        );

    \I__6820\ : Span4Mux_v
    port map (
            O => \N__34825\,
            I => \N__34817\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__34822\,
            I => \N__34817\
        );

    \I__6818\ : Odrv4
    port map (
            O => \N__34817\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__6817\ : InMux
    port map (
            O => \N__34814\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__6816\ : CascadeMux
    port map (
            O => \N__34811\,
            I => \N__34808\
        );

    \I__6815\ : InMux
    port map (
            O => \N__34808\,
            I => \N__34804\
        );

    \I__6814\ : InMux
    port map (
            O => \N__34807\,
            I => \N__34801\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__34804\,
            I => \N__34795\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__34801\,
            I => \N__34795\
        );

    \I__6811\ : InMux
    port map (
            O => \N__34800\,
            I => \N__34792\
        );

    \I__6810\ : Span4Mux_h
    port map (
            O => \N__34795\,
            I => \N__34789\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__34792\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__6808\ : Odrv4
    port map (
            O => \N__34789\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__6807\ : InMux
    port map (
            O => \N__34784\,
            I => \N__34781\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__34781\,
            I => \N__34778\
        );

    \I__6805\ : Span4Mux_v
    port map (
            O => \N__34778\,
            I => \N__34773\
        );

    \I__6804\ : InMux
    port map (
            O => \N__34777\,
            I => \N__34770\
        );

    \I__6803\ : InMux
    port map (
            O => \N__34776\,
            I => \N__34767\
        );

    \I__6802\ : Span4Mux_v
    port map (
            O => \N__34773\,
            I => \N__34759\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__34770\,
            I => \N__34759\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__34767\,
            I => \N__34759\
        );

    \I__6799\ : InMux
    port map (
            O => \N__34766\,
            I => \N__34756\
        );

    \I__6798\ : Span4Mux_h
    port map (
            O => \N__34759\,
            I => \N__34751\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__34756\,
            I => \N__34751\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__34751\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__6795\ : InMux
    port map (
            O => \N__34748\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__6794\ : CascadeMux
    port map (
            O => \N__34745\,
            I => \N__34742\
        );

    \I__6793\ : InMux
    port map (
            O => \N__34742\,
            I => \N__34738\
        );

    \I__6792\ : InMux
    port map (
            O => \N__34741\,
            I => \N__34735\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__34738\,
            I => \N__34729\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__34735\,
            I => \N__34729\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34726\
        );

    \I__6788\ : Span4Mux_h
    port map (
            O => \N__34729\,
            I => \N__34723\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__34726\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__6786\ : Odrv4
    port map (
            O => \N__34723\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34718\,
            I => \N__34713\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34717\,
            I => \N__34710\
        );

    \I__6783\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34707\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__34713\,
            I => \N__34703\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__34710\,
            I => \N__34698\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__34707\,
            I => \N__34698\
        );

    \I__6779\ : InMux
    port map (
            O => \N__34706\,
            I => \N__34695\
        );

    \I__6778\ : Span4Mux_v
    port map (
            O => \N__34703\,
            I => \N__34690\
        );

    \I__6777\ : Span4Mux_v
    port map (
            O => \N__34698\,
            I => \N__34690\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__34695\,
            I => \N__34687\
        );

    \I__6775\ : Span4Mux_h
    port map (
            O => \N__34690\,
            I => \N__34684\
        );

    \I__6774\ : Span4Mux_v
    port map (
            O => \N__34687\,
            I => \N__34681\
        );

    \I__6773\ : Odrv4
    port map (
            O => \N__34684\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__6772\ : Odrv4
    port map (
            O => \N__34681\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__6771\ : InMux
    port map (
            O => \N__34676\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__6770\ : CascadeMux
    port map (
            O => \N__34673\,
            I => \N__34670\
        );

    \I__6769\ : InMux
    port map (
            O => \N__34670\,
            I => \N__34666\
        );

    \I__6768\ : InMux
    port map (
            O => \N__34669\,
            I => \N__34663\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__34666\,
            I => \N__34657\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__34663\,
            I => \N__34657\
        );

    \I__6765\ : InMux
    port map (
            O => \N__34662\,
            I => \N__34654\
        );

    \I__6764\ : Span4Mux_h
    port map (
            O => \N__34657\,
            I => \N__34651\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__34654\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__6762\ : Odrv4
    port map (
            O => \N__34651\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__6761\ : InMux
    port map (
            O => \N__34646\,
            I => \N__34641\
        );

    \I__6760\ : InMux
    port map (
            O => \N__34645\,
            I => \N__34637\
        );

    \I__6759\ : CascadeMux
    port map (
            O => \N__34644\,
            I => \N__34634\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__34641\,
            I => \N__34631\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34640\,
            I => \N__34628\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__34637\,
            I => \N__34625\
        );

    \I__6755\ : InMux
    port map (
            O => \N__34634\,
            I => \N__34622\
        );

    \I__6754\ : Span4Mux_h
    port map (
            O => \N__34631\,
            I => \N__34617\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__34628\,
            I => \N__34617\
        );

    \I__6752\ : Span4Mux_h
    port map (
            O => \N__34625\,
            I => \N__34612\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__34622\,
            I => \N__34612\
        );

    \I__6750\ : Span4Mux_h
    port map (
            O => \N__34617\,
            I => \N__34609\
        );

    \I__6749\ : Span4Mux_v
    port map (
            O => \N__34612\,
            I => \N__34606\
        );

    \I__6748\ : Odrv4
    port map (
            O => \N__34609\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__6747\ : Odrv4
    port map (
            O => \N__34606\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__6746\ : InMux
    port map (
            O => \N__34601\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__6745\ : InMux
    port map (
            O => \N__34598\,
            I => \N__34592\
        );

    \I__6744\ : InMux
    port map (
            O => \N__34597\,
            I => \N__34592\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__34592\,
            I => \N__34588\
        );

    \I__6742\ : InMux
    port map (
            O => \N__34591\,
            I => \N__34585\
        );

    \I__6741\ : Span4Mux_h
    port map (
            O => \N__34588\,
            I => \N__34582\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__34585\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__6739\ : Odrv4
    port map (
            O => \N__34582\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__6738\ : InMux
    port map (
            O => \N__34577\,
            I => \N__34573\
        );

    \I__6737\ : InMux
    port map (
            O => \N__34576\,
            I => \N__34570\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__34573\,
            I => \N__34567\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__34570\,
            I => \N__34562\
        );

    \I__6734\ : Span4Mux_v
    port map (
            O => \N__34567\,
            I => \N__34559\
        );

    \I__6733\ : InMux
    port map (
            O => \N__34566\,
            I => \N__34556\
        );

    \I__6732\ : InMux
    port map (
            O => \N__34565\,
            I => \N__34553\
        );

    \I__6731\ : Span4Mux_h
    port map (
            O => \N__34562\,
            I => \N__34546\
        );

    \I__6730\ : Span4Mux_h
    port map (
            O => \N__34559\,
            I => \N__34546\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__34556\,
            I => \N__34546\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__34553\,
            I => \N__34543\
        );

    \I__6727\ : Odrv4
    port map (
            O => \N__34546\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__6726\ : Odrv4
    port map (
            O => \N__34543\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__6725\ : InMux
    port map (
            O => \N__34538\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__6724\ : InMux
    port map (
            O => \N__34535\,
            I => \N__34529\
        );

    \I__6723\ : InMux
    port map (
            O => \N__34534\,
            I => \N__34529\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__34529\,
            I => \N__34525\
        );

    \I__6721\ : InMux
    port map (
            O => \N__34528\,
            I => \N__34522\
        );

    \I__6720\ : Span4Mux_h
    port map (
            O => \N__34525\,
            I => \N__34519\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__34522\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__6718\ : Odrv4
    port map (
            O => \N__34519\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__6717\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34509\
        );

    \I__6716\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34505\
        );

    \I__6715\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34502\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__34509\,
            I => \N__34499\
        );

    \I__6713\ : InMux
    port map (
            O => \N__34508\,
            I => \N__34496\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34493\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__34502\,
            I => \N__34490\
        );

    \I__6710\ : Span4Mux_v
    port map (
            O => \N__34499\,
            I => \N__34485\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__34496\,
            I => \N__34485\
        );

    \I__6708\ : Span4Mux_h
    port map (
            O => \N__34493\,
            I => \N__34482\
        );

    \I__6707\ : Span4Mux_h
    port map (
            O => \N__34490\,
            I => \N__34479\
        );

    \I__6706\ : Odrv4
    port map (
            O => \N__34485\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__6705\ : Odrv4
    port map (
            O => \N__34482\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__6704\ : Odrv4
    port map (
            O => \N__34479\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__6703\ : InMux
    port map (
            O => \N__34472\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__6702\ : InMux
    port map (
            O => \N__34469\,
            I => \N__34464\
        );

    \I__6701\ : InMux
    port map (
            O => \N__34468\,
            I => \N__34459\
        );

    \I__6700\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34459\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__34464\,
            I => \N__34453\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__34459\,
            I => \N__34453\
        );

    \I__6697\ : InMux
    port map (
            O => \N__34458\,
            I => \N__34450\
        );

    \I__6696\ : Span4Mux_v
    port map (
            O => \N__34453\,
            I => \N__34445\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__34450\,
            I => \N__34445\
        );

    \I__6694\ : Span4Mux_h
    port map (
            O => \N__34445\,
            I => \N__34442\
        );

    \I__6693\ : Odrv4
    port map (
            O => \N__34442\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__6692\ : InMux
    port map (
            O => \N__34439\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__6691\ : CascadeMux
    port map (
            O => \N__34436\,
            I => \N__34433\
        );

    \I__6690\ : InMux
    port map (
            O => \N__34433\,
            I => \N__34430\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__34430\,
            I => \N__34425\
        );

    \I__6688\ : InMux
    port map (
            O => \N__34429\,
            I => \N__34422\
        );

    \I__6687\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34419\
        );

    \I__6686\ : Span4Mux_v
    port map (
            O => \N__34425\,
            I => \N__34416\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__34422\,
            I => \N__34413\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__34419\,
            I => \N__34408\
        );

    \I__6683\ : Span4Mux_h
    port map (
            O => \N__34416\,
            I => \N__34408\
        );

    \I__6682\ : Span4Mux_h
    port map (
            O => \N__34413\,
            I => \N__34405\
        );

    \I__6681\ : Odrv4
    port map (
            O => \N__34408\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__6680\ : Odrv4
    port map (
            O => \N__34405\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__6679\ : CascadeMux
    port map (
            O => \N__34400\,
            I => \N__34397\
        );

    \I__6678\ : InMux
    port map (
            O => \N__34397\,
            I => \N__34392\
        );

    \I__6677\ : InMux
    port map (
            O => \N__34396\,
            I => \N__34389\
        );

    \I__6676\ : InMux
    port map (
            O => \N__34395\,
            I => \N__34386\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__34392\,
            I => \N__34380\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__34389\,
            I => \N__34380\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__34386\,
            I => \N__34377\
        );

    \I__6672\ : InMux
    port map (
            O => \N__34385\,
            I => \N__34374\
        );

    \I__6671\ : Span4Mux_v
    port map (
            O => \N__34380\,
            I => \N__34371\
        );

    \I__6670\ : Span4Mux_h
    port map (
            O => \N__34377\,
            I => \N__34366\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__34374\,
            I => \N__34366\
        );

    \I__6668\ : Span4Mux_h
    port map (
            O => \N__34371\,
            I => \N__34363\
        );

    \I__6667\ : Span4Mux_v
    port map (
            O => \N__34366\,
            I => \N__34360\
        );

    \I__6666\ : Odrv4
    port map (
            O => \N__34363\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__6665\ : Odrv4
    port map (
            O => \N__34360\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__6664\ : InMux
    port map (
            O => \N__34355\,
            I => \bfn_13_11_0_\
        );

    \I__6663\ : CascadeMux
    port map (
            O => \N__34352\,
            I => \N__34349\
        );

    \I__6662\ : InMux
    port map (
            O => \N__34349\,
            I => \N__34344\
        );

    \I__6661\ : InMux
    port map (
            O => \N__34348\,
            I => \N__34341\
        );

    \I__6660\ : InMux
    port map (
            O => \N__34347\,
            I => \N__34338\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__34344\,
            I => \N__34335\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__34341\,
            I => \N__34332\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__34338\,
            I => \N__34327\
        );

    \I__6656\ : Span4Mux_v
    port map (
            O => \N__34335\,
            I => \N__34327\
        );

    \I__6655\ : Span4Mux_h
    port map (
            O => \N__34332\,
            I => \N__34324\
        );

    \I__6654\ : Odrv4
    port map (
            O => \N__34327\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__6653\ : Odrv4
    port map (
            O => \N__34324\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__6652\ : CascadeMux
    port map (
            O => \N__34319\,
            I => \N__34316\
        );

    \I__6651\ : InMux
    port map (
            O => \N__34316\,
            I => \N__34311\
        );

    \I__6650\ : InMux
    port map (
            O => \N__34315\,
            I => \N__34308\
        );

    \I__6649\ : CascadeMux
    port map (
            O => \N__34314\,
            I => \N__34305\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__34311\,
            I => \N__34301\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__34308\,
            I => \N__34298\
        );

    \I__6646\ : InMux
    port map (
            O => \N__34305\,
            I => \N__34295\
        );

    \I__6645\ : InMux
    port map (
            O => \N__34304\,
            I => \N__34292\
        );

    \I__6644\ : Span4Mux_v
    port map (
            O => \N__34301\,
            I => \N__34285\
        );

    \I__6643\ : Span4Mux_h
    port map (
            O => \N__34298\,
            I => \N__34285\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__34295\,
            I => \N__34285\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__34292\,
            I => \N__34282\
        );

    \I__6640\ : Span4Mux_h
    port map (
            O => \N__34285\,
            I => \N__34279\
        );

    \I__6639\ : Odrv12
    port map (
            O => \N__34282\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__6638\ : Odrv4
    port map (
            O => \N__34279\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__6637\ : InMux
    port map (
            O => \N__34274\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__6636\ : CascadeMux
    port map (
            O => \N__34271\,
            I => \N__34268\
        );

    \I__6635\ : InMux
    port map (
            O => \N__34268\,
            I => \N__34264\
        );

    \I__6634\ : InMux
    port map (
            O => \N__34267\,
            I => \N__34261\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__34264\,
            I => \N__34255\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__34261\,
            I => \N__34255\
        );

    \I__6631\ : InMux
    port map (
            O => \N__34260\,
            I => \N__34252\
        );

    \I__6630\ : Span4Mux_h
    port map (
            O => \N__34255\,
            I => \N__34249\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__34252\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__34249\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__6627\ : InMux
    port map (
            O => \N__34244\,
            I => \N__34240\
        );

    \I__6626\ : InMux
    port map (
            O => \N__34243\,
            I => \N__34236\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__34240\,
            I => \N__34233\
        );

    \I__6624\ : InMux
    port map (
            O => \N__34239\,
            I => \N__34230\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__34236\,
            I => \N__34226\
        );

    \I__6622\ : Span4Mux_v
    port map (
            O => \N__34233\,
            I => \N__34221\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__34230\,
            I => \N__34221\
        );

    \I__6620\ : InMux
    port map (
            O => \N__34229\,
            I => \N__34218\
        );

    \I__6619\ : Span4Mux_v
    port map (
            O => \N__34226\,
            I => \N__34215\
        );

    \I__6618\ : Span4Mux_h
    port map (
            O => \N__34221\,
            I => \N__34210\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__34218\,
            I => \N__34210\
        );

    \I__6616\ : Odrv4
    port map (
            O => \N__34215\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__6615\ : Odrv4
    port map (
            O => \N__34210\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__6614\ : InMux
    port map (
            O => \N__34205\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__6613\ : CascadeMux
    port map (
            O => \N__34202\,
            I => \N__34199\
        );

    \I__6612\ : InMux
    port map (
            O => \N__34199\,
            I => \N__34195\
        );

    \I__6611\ : InMux
    port map (
            O => \N__34198\,
            I => \N__34192\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__34195\,
            I => \N__34186\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__34192\,
            I => \N__34186\
        );

    \I__6608\ : InMux
    port map (
            O => \N__34191\,
            I => \N__34183\
        );

    \I__6607\ : Span4Mux_h
    port map (
            O => \N__34186\,
            I => \N__34180\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__34183\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__6605\ : Odrv4
    port map (
            O => \N__34180\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__6604\ : InMux
    port map (
            O => \N__34175\,
            I => \N__34170\
        );

    \I__6603\ : InMux
    port map (
            O => \N__34174\,
            I => \N__34167\
        );

    \I__6602\ : CascadeMux
    port map (
            O => \N__34173\,
            I => \N__34163\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__34170\,
            I => \N__34160\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__34167\,
            I => \N__34157\
        );

    \I__6599\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34154\
        );

    \I__6598\ : InMux
    port map (
            O => \N__34163\,
            I => \N__34151\
        );

    \I__6597\ : Span4Mux_h
    port map (
            O => \N__34160\,
            I => \N__34144\
        );

    \I__6596\ : Span4Mux_h
    port map (
            O => \N__34157\,
            I => \N__34144\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__34154\,
            I => \N__34144\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__34151\,
            I => \N__34141\
        );

    \I__6593\ : Odrv4
    port map (
            O => \N__34144\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__6592\ : Odrv4
    port map (
            O => \N__34141\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__6591\ : InMux
    port map (
            O => \N__34136\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__6590\ : CascadeMux
    port map (
            O => \N__34133\,
            I => \N__34130\
        );

    \I__6589\ : InMux
    port map (
            O => \N__34130\,
            I => \N__34126\
        );

    \I__6588\ : InMux
    port map (
            O => \N__34129\,
            I => \N__34123\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__34126\,
            I => \N__34117\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__34123\,
            I => \N__34117\
        );

    \I__6585\ : InMux
    port map (
            O => \N__34122\,
            I => \N__34114\
        );

    \I__6584\ : Span4Mux_h
    port map (
            O => \N__34117\,
            I => \N__34111\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__34114\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__6582\ : Odrv4
    port map (
            O => \N__34111\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__6581\ : InMux
    port map (
            O => \N__34106\,
            I => \N__34103\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__34103\,
            I => \N__34097\
        );

    \I__6579\ : InMux
    port map (
            O => \N__34102\,
            I => \N__34092\
        );

    \I__6578\ : InMux
    port map (
            O => \N__34101\,
            I => \N__34092\
        );

    \I__6577\ : InMux
    port map (
            O => \N__34100\,
            I => \N__34089\
        );

    \I__6576\ : Span4Mux_v
    port map (
            O => \N__34097\,
            I => \N__34082\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__34092\,
            I => \N__34082\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__34089\,
            I => \N__34082\
        );

    \I__6573\ : Span4Mux_h
    port map (
            O => \N__34082\,
            I => \N__34079\
        );

    \I__6572\ : Odrv4
    port map (
            O => \N__34079\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__6571\ : InMux
    port map (
            O => \N__34076\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__6570\ : CascadeMux
    port map (
            O => \N__34073\,
            I => \N__34070\
        );

    \I__6569\ : InMux
    port map (
            O => \N__34070\,
            I => \N__34066\
        );

    \I__6568\ : InMux
    port map (
            O => \N__34069\,
            I => \N__34063\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__34066\,
            I => \N__34057\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__34063\,
            I => \N__34057\
        );

    \I__6565\ : InMux
    port map (
            O => \N__34062\,
            I => \N__34054\
        );

    \I__6564\ : Span4Mux_h
    port map (
            O => \N__34057\,
            I => \N__34051\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__34054\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__34051\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__6561\ : InMux
    port map (
            O => \N__34046\,
            I => \N__34041\
        );

    \I__6560\ : InMux
    port map (
            O => \N__34045\,
            I => \N__34038\
        );

    \I__6559\ : InMux
    port map (
            O => \N__34044\,
            I => \N__34035\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__34041\,
            I => \N__34030\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__34038\,
            I => \N__34030\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__34035\,
            I => \N__34026\
        );

    \I__6555\ : Span4Mux_v
    port map (
            O => \N__34030\,
            I => \N__34023\
        );

    \I__6554\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34020\
        );

    \I__6553\ : Span4Mux_h
    port map (
            O => \N__34026\,
            I => \N__34017\
        );

    \I__6552\ : Sp12to4
    port map (
            O => \N__34023\,
            I => \N__34014\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__34020\,
            I => \N__34011\
        );

    \I__6550\ : Odrv4
    port map (
            O => \N__34017\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__6549\ : Odrv12
    port map (
            O => \N__34014\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__6548\ : Odrv4
    port map (
            O => \N__34011\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__6547\ : InMux
    port map (
            O => \N__34004\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__6546\ : CascadeMux
    port map (
            O => \N__34001\,
            I => \N__33998\
        );

    \I__6545\ : InMux
    port map (
            O => \N__33998\,
            I => \N__33994\
        );

    \I__6544\ : InMux
    port map (
            O => \N__33997\,
            I => \N__33991\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__33994\,
            I => \N__33985\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__33991\,
            I => \N__33985\
        );

    \I__6541\ : InMux
    port map (
            O => \N__33990\,
            I => \N__33982\
        );

    \I__6540\ : Span4Mux_h
    port map (
            O => \N__33985\,
            I => \N__33979\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__33982\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__6538\ : Odrv4
    port map (
            O => \N__33979\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__6537\ : InMux
    port map (
            O => \N__33974\,
            I => \N__33971\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__33971\,
            I => \N__33966\
        );

    \I__6535\ : InMux
    port map (
            O => \N__33970\,
            I => \N__33961\
        );

    \I__6534\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33961\
        );

    \I__6533\ : Span4Mux_v
    port map (
            O => \N__33966\,
            I => \N__33955\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__33961\,
            I => \N__33955\
        );

    \I__6531\ : InMux
    port map (
            O => \N__33960\,
            I => \N__33952\
        );

    \I__6530\ : Span4Mux_h
    port map (
            O => \N__33955\,
            I => \N__33947\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__33952\,
            I => \N__33947\
        );

    \I__6528\ : Sp12to4
    port map (
            O => \N__33947\,
            I => \N__33944\
        );

    \I__6527\ : Odrv12
    port map (
            O => \N__33944\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__6526\ : InMux
    port map (
            O => \N__33941\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__6525\ : CascadeMux
    port map (
            O => \N__33938\,
            I => \N__33935\
        );

    \I__6524\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33931\
        );

    \I__6523\ : InMux
    port map (
            O => \N__33934\,
            I => \N__33928\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__33931\,
            I => \N__33924\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__33928\,
            I => \N__33921\
        );

    \I__6520\ : InMux
    port map (
            O => \N__33927\,
            I => \N__33918\
        );

    \I__6519\ : Span4Mux_v
    port map (
            O => \N__33924\,
            I => \N__33915\
        );

    \I__6518\ : Odrv12
    port map (
            O => \N__33921\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__33918\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__6516\ : Odrv4
    port map (
            O => \N__33915\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__6515\ : InMux
    port map (
            O => \N__33908\,
            I => \N__33904\
        );

    \I__6514\ : InMux
    port map (
            O => \N__33907\,
            I => \N__33899\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__33904\,
            I => \N__33896\
        );

    \I__6512\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33891\
        );

    \I__6511\ : InMux
    port map (
            O => \N__33902\,
            I => \N__33891\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33888\
        );

    \I__6509\ : Span4Mux_v
    port map (
            O => \N__33896\,
            I => \N__33885\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__33891\,
            I => \N__33882\
        );

    \I__6507\ : Span4Mux_h
    port map (
            O => \N__33888\,
            I => \N__33879\
        );

    \I__6506\ : Sp12to4
    port map (
            O => \N__33885\,
            I => \N__33874\
        );

    \I__6505\ : Span12Mux_s9_v
    port map (
            O => \N__33882\,
            I => \N__33874\
        );

    \I__6504\ : Odrv4
    port map (
            O => \N__33879\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__6503\ : Odrv12
    port map (
            O => \N__33874\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__6502\ : CascadeMux
    port map (
            O => \N__33869\,
            I => \N__33866\
        );

    \I__6501\ : InMux
    port map (
            O => \N__33866\,
            I => \N__33861\
        );

    \I__6500\ : InMux
    port map (
            O => \N__33865\,
            I => \N__33858\
        );

    \I__6499\ : InMux
    port map (
            O => \N__33864\,
            I => \N__33855\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__33861\,
            I => \N__33852\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__33858\,
            I => \N__33849\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__33855\,
            I => \N__33844\
        );

    \I__6495\ : Span4Mux_v
    port map (
            O => \N__33852\,
            I => \N__33844\
        );

    \I__6494\ : Odrv12
    port map (
            O => \N__33849\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__6493\ : Odrv4
    port map (
            O => \N__33844\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__6492\ : CascadeMux
    port map (
            O => \N__33839\,
            I => \N__33835\
        );

    \I__6491\ : InMux
    port map (
            O => \N__33838\,
            I => \N__33831\
        );

    \I__6490\ : InMux
    port map (
            O => \N__33835\,
            I => \N__33827\
        );

    \I__6489\ : InMux
    port map (
            O => \N__33834\,
            I => \N__33824\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__33831\,
            I => \N__33821\
        );

    \I__6487\ : InMux
    port map (
            O => \N__33830\,
            I => \N__33818\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__33827\,
            I => \N__33815\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__33824\,
            I => \N__33808\
        );

    \I__6484\ : Span4Mux_h
    port map (
            O => \N__33821\,
            I => \N__33808\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__33818\,
            I => \N__33808\
        );

    \I__6482\ : Span4Mux_h
    port map (
            O => \N__33815\,
            I => \N__33805\
        );

    \I__6481\ : Span4Mux_h
    port map (
            O => \N__33808\,
            I => \N__33802\
        );

    \I__6480\ : Span4Mux_h
    port map (
            O => \N__33805\,
            I => \N__33799\
        );

    \I__6479\ : Odrv4
    port map (
            O => \N__33802\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__6478\ : Odrv4
    port map (
            O => \N__33799\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__6477\ : InMux
    port map (
            O => \N__33794\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__6476\ : InMux
    port map (
            O => \N__33791\,
            I => \N__33785\
        );

    \I__6475\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33785\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__33785\,
            I => \N__33781\
        );

    \I__6473\ : InMux
    port map (
            O => \N__33784\,
            I => \N__33778\
        );

    \I__6472\ : Span4Mux_h
    port map (
            O => \N__33781\,
            I => \N__33775\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__33778\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__6470\ : Odrv4
    port map (
            O => \N__33775\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__6469\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33765\
        );

    \I__6468\ : InMux
    port map (
            O => \N__33769\,
            I => \N__33762\
        );

    \I__6467\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33759\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__33765\,
            I => \N__33755\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__33762\,
            I => \N__33752\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__33759\,
            I => \N__33749\
        );

    \I__6463\ : InMux
    port map (
            O => \N__33758\,
            I => \N__33746\
        );

    \I__6462\ : Span4Mux_v
    port map (
            O => \N__33755\,
            I => \N__33743\
        );

    \I__6461\ : Span4Mux_h
    port map (
            O => \N__33752\,
            I => \N__33740\
        );

    \I__6460\ : Span4Mux_v
    port map (
            O => \N__33749\,
            I => \N__33737\
        );

    \I__6459\ : LocalMux
    port map (
            O => \N__33746\,
            I => \N__33734\
        );

    \I__6458\ : Span4Mux_h
    port map (
            O => \N__33743\,
            I => \N__33729\
        );

    \I__6457\ : Span4Mux_v
    port map (
            O => \N__33740\,
            I => \N__33729\
        );

    \I__6456\ : Span4Mux_h
    port map (
            O => \N__33737\,
            I => \N__33724\
        );

    \I__6455\ : Span4Mux_v
    port map (
            O => \N__33734\,
            I => \N__33724\
        );

    \I__6454\ : Odrv4
    port map (
            O => \N__33729\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__6453\ : Odrv4
    port map (
            O => \N__33724\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__6452\ : InMux
    port map (
            O => \N__33719\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__33716\,
            I => \N__33713\
        );

    \I__6450\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33709\
        );

    \I__6449\ : InMux
    port map (
            O => \N__33712\,
            I => \N__33706\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__33709\,
            I => \N__33700\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__33706\,
            I => \N__33700\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33705\,
            I => \N__33697\
        );

    \I__6445\ : Span4Mux_h
    port map (
            O => \N__33700\,
            I => \N__33694\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__33697\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__6443\ : Odrv4
    port map (
            O => \N__33694\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__6442\ : InMux
    port map (
            O => \N__33689\,
            I => \N__33684\
        );

    \I__6441\ : InMux
    port map (
            O => \N__33688\,
            I => \N__33680\
        );

    \I__6440\ : InMux
    port map (
            O => \N__33687\,
            I => \N__33677\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__33684\,
            I => \N__33674\
        );

    \I__6438\ : InMux
    port map (
            O => \N__33683\,
            I => \N__33671\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__33680\,
            I => \N__33666\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__33677\,
            I => \N__33666\
        );

    \I__6435\ : Span4Mux_v
    port map (
            O => \N__33674\,
            I => \N__33663\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__33671\,
            I => \N__33660\
        );

    \I__6433\ : Span4Mux_v
    port map (
            O => \N__33666\,
            I => \N__33657\
        );

    \I__6432\ : Span4Mux_h
    port map (
            O => \N__33663\,
            I => \N__33652\
        );

    \I__6431\ : Span4Mux_v
    port map (
            O => \N__33660\,
            I => \N__33652\
        );

    \I__6430\ : Odrv4
    port map (
            O => \N__33657\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__6429\ : Odrv4
    port map (
            O => \N__33652\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__6428\ : InMux
    port map (
            O => \N__33647\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__6427\ : CascadeMux
    port map (
            O => \N__33644\,
            I => \N__33640\
        );

    \I__6426\ : InMux
    port map (
            O => \N__33643\,
            I => \N__33637\
        );

    \I__6425\ : InMux
    port map (
            O => \N__33640\,
            I => \N__33634\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__33637\,
            I => \N__33628\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__33634\,
            I => \N__33628\
        );

    \I__6422\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33625\
        );

    \I__6421\ : Span4Mux_h
    port map (
            O => \N__33628\,
            I => \N__33622\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__33625\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__6419\ : Odrv4
    port map (
            O => \N__33622\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__6418\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33613\
        );

    \I__6417\ : InMux
    port map (
            O => \N__33616\,
            I => \N__33610\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__33613\,
            I => \N__33603\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__33610\,
            I => \N__33603\
        );

    \I__6414\ : InMux
    port map (
            O => \N__33609\,
            I => \N__33600\
        );

    \I__6413\ : InMux
    port map (
            O => \N__33608\,
            I => \N__33597\
        );

    \I__6412\ : Span4Mux_v
    port map (
            O => \N__33603\,
            I => \N__33594\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__33600\,
            I => \N__33591\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__33597\,
            I => \N__33588\
        );

    \I__6409\ : Span4Mux_h
    port map (
            O => \N__33594\,
            I => \N__33585\
        );

    \I__6408\ : Span4Mux_v
    port map (
            O => \N__33591\,
            I => \N__33580\
        );

    \I__6407\ : Span4Mux_v
    port map (
            O => \N__33588\,
            I => \N__33580\
        );

    \I__6406\ : Odrv4
    port map (
            O => \N__33585\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__6405\ : Odrv4
    port map (
            O => \N__33580\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__6404\ : InMux
    port map (
            O => \N__33575\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__6403\ : CascadeMux
    port map (
            O => \N__33572\,
            I => \N__33569\
        );

    \I__6402\ : InMux
    port map (
            O => \N__33569\,
            I => \N__33565\
        );

    \I__6401\ : InMux
    port map (
            O => \N__33568\,
            I => \N__33562\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__33565\,
            I => \N__33556\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__33562\,
            I => \N__33556\
        );

    \I__6398\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33553\
        );

    \I__6397\ : Span4Mux_h
    port map (
            O => \N__33556\,
            I => \N__33550\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__33553\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__6395\ : Odrv4
    port map (
            O => \N__33550\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__6394\ : InMux
    port map (
            O => \N__33545\,
            I => \N__33539\
        );

    \I__6393\ : InMux
    port map (
            O => \N__33544\,
            I => \N__33539\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__33539\,
            I => \N__33534\
        );

    \I__6391\ : InMux
    port map (
            O => \N__33538\,
            I => \N__33531\
        );

    \I__6390\ : InMux
    port map (
            O => \N__33537\,
            I => \N__33528\
        );

    \I__6389\ : Span4Mux_h
    port map (
            O => \N__33534\,
            I => \N__33525\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__33531\,
            I => \N__33522\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__33528\,
            I => \N__33519\
        );

    \I__6386\ : Span4Mux_h
    port map (
            O => \N__33525\,
            I => \N__33516\
        );

    \I__6385\ : Span4Mux_h
    port map (
            O => \N__33522\,
            I => \N__33511\
        );

    \I__6384\ : Span4Mux_h
    port map (
            O => \N__33519\,
            I => \N__33511\
        );

    \I__6383\ : Odrv4
    port map (
            O => \N__33516\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__6382\ : Odrv4
    port map (
            O => \N__33511\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__6381\ : InMux
    port map (
            O => \N__33506\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__6380\ : CascadeMux
    port map (
            O => \N__33503\,
            I => \N__33499\
        );

    \I__6379\ : CascadeMux
    port map (
            O => \N__33502\,
            I => \N__33496\
        );

    \I__6378\ : InMux
    port map (
            O => \N__33499\,
            I => \N__33491\
        );

    \I__6377\ : InMux
    port map (
            O => \N__33496\,
            I => \N__33491\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__33491\,
            I => \N__33487\
        );

    \I__6375\ : InMux
    port map (
            O => \N__33490\,
            I => \N__33484\
        );

    \I__6374\ : Span4Mux_h
    port map (
            O => \N__33487\,
            I => \N__33481\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__33484\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__6372\ : Odrv4
    port map (
            O => \N__33481\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__6371\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33471\
        );

    \I__6370\ : InMux
    port map (
            O => \N__33475\,
            I => \N__33466\
        );

    \I__6369\ : InMux
    port map (
            O => \N__33474\,
            I => \N__33466\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__33471\,
            I => \N__33462\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__33466\,
            I => \N__33459\
        );

    \I__6366\ : InMux
    port map (
            O => \N__33465\,
            I => \N__33456\
        );

    \I__6365\ : Span4Mux_v
    port map (
            O => \N__33462\,
            I => \N__33453\
        );

    \I__6364\ : Span4Mux_h
    port map (
            O => \N__33459\,
            I => \N__33450\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__33456\,
            I => \N__33447\
        );

    \I__6362\ : Span4Mux_h
    port map (
            O => \N__33453\,
            I => \N__33444\
        );

    \I__6361\ : Span4Mux_h
    port map (
            O => \N__33450\,
            I => \N__33441\
        );

    \I__6360\ : Span4Mux_v
    port map (
            O => \N__33447\,
            I => \N__33438\
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__33444\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__6358\ : Odrv4
    port map (
            O => \N__33441\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__6357\ : Odrv4
    port map (
            O => \N__33438\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__6356\ : InMux
    port map (
            O => \N__33431\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__6355\ : CascadeMux
    port map (
            O => \N__33428\,
            I => \N__33425\
        );

    \I__6354\ : InMux
    port map (
            O => \N__33425\,
            I => \N__33421\
        );

    \I__6353\ : InMux
    port map (
            O => \N__33424\,
            I => \N__33418\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__33421\,
            I => \N__33412\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__33418\,
            I => \N__33412\
        );

    \I__6350\ : InMux
    port map (
            O => \N__33417\,
            I => \N__33409\
        );

    \I__6349\ : Span4Mux_h
    port map (
            O => \N__33412\,
            I => \N__33406\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__33409\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__6347\ : Odrv4
    port map (
            O => \N__33406\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__6346\ : CascadeMux
    port map (
            O => \N__33401\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5_cascade_\
        );

    \I__6345\ : CascadeMux
    port map (
            O => \N__33398\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\
        );

    \I__6344\ : InMux
    port map (
            O => \N__33395\,
            I => \N__33392\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__33392\,
            I => \N__33389\
        );

    \I__6342\ : Odrv12
    port map (
            O => \N__33389\,
            I => \phase_controller_inst1.test_0_sqmuxa\
        );

    \I__6341\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33380\
        );

    \I__6340\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33380\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__33380\,
            I => \N__33377\
        );

    \I__6338\ : Odrv4
    port map (
            O => \N__33377\,
            I => \phase_controller_inst1.N_56\
        );

    \I__6337\ : CascadeMux
    port map (
            O => \N__33374\,
            I => \N__33371\
        );

    \I__6336\ : InMux
    port map (
            O => \N__33371\,
            I => \N__33367\
        );

    \I__6335\ : InMux
    port map (
            O => \N__33370\,
            I => \N__33364\
        );

    \I__6334\ : LocalMux
    port map (
            O => \N__33367\,
            I => \N__33360\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__33364\,
            I => \N__33357\
        );

    \I__6332\ : InMux
    port map (
            O => \N__33363\,
            I => \N__33354\
        );

    \I__6331\ : Span4Mux_h
    port map (
            O => \N__33360\,
            I => \N__33348\
        );

    \I__6330\ : Span12Mux_h
    port map (
            O => \N__33357\,
            I => \N__33345\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__33354\,
            I => \N__33342\
        );

    \I__6328\ : InMux
    port map (
            O => \N__33353\,
            I => \N__33337\
        );

    \I__6327\ : InMux
    port map (
            O => \N__33352\,
            I => \N__33337\
        );

    \I__6326\ : InMux
    port map (
            O => \N__33351\,
            I => \N__33334\
        );

    \I__6325\ : Span4Mux_v
    port map (
            O => \N__33348\,
            I => \N__33331\
        );

    \I__6324\ : Span12Mux_v
    port map (
            O => \N__33345\,
            I => \N__33328\
        );

    \I__6323\ : Span4Mux_h
    port map (
            O => \N__33342\,
            I => \N__33325\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__33337\,
            I => phase_controller_inst1_state_4
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__33334\,
            I => phase_controller_inst1_state_4
        );

    \I__6320\ : Odrv4
    port map (
            O => \N__33331\,
            I => phase_controller_inst1_state_4
        );

    \I__6319\ : Odrv12
    port map (
            O => \N__33328\,
            I => phase_controller_inst1_state_4
        );

    \I__6318\ : Odrv4
    port map (
            O => \N__33325\,
            I => phase_controller_inst1_state_4
        );

    \I__6317\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33311\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__33311\,
            I => \N__33308\
        );

    \I__6315\ : Odrv4
    port map (
            O => \N__33308\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\
        );

    \I__6314\ : InMux
    port map (
            O => \N__33305\,
            I => \current_shift_inst.control_input_cry_24\
        );

    \I__6313\ : CascadeMux
    port map (
            O => \N__33302\,
            I => \N__33299\
        );

    \I__6312\ : InMux
    port map (
            O => \N__33299\,
            I => \N__33296\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__33296\,
            I => \N__33293\
        );

    \I__6310\ : Odrv4
    port map (
            O => \N__33293\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\
        );

    \I__6309\ : InMux
    port map (
            O => \N__33290\,
            I => \current_shift_inst.control_input_cry_25\
        );

    \I__6308\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33284\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__33284\,
            I => \N__33281\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__33281\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\
        );

    \I__6305\ : InMux
    port map (
            O => \N__33278\,
            I => \current_shift_inst.control_input_cry_26\
        );

    \I__6304\ : InMux
    port map (
            O => \N__33275\,
            I => \N__33272\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__33272\,
            I => \N__33269\
        );

    \I__6302\ : Odrv4
    port map (
            O => \N__33269\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\
        );

    \I__6301\ : InMux
    port map (
            O => \N__33266\,
            I => \current_shift_inst.control_input_cry_27\
        );

    \I__6300\ : CascadeMux
    port map (
            O => \N__33263\,
            I => \N__33260\
        );

    \I__6299\ : InMux
    port map (
            O => \N__33260\,
            I => \N__33257\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__33257\,
            I => \N__33254\
        );

    \I__6297\ : Odrv4
    port map (
            O => \N__33254\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\
        );

    \I__6296\ : InMux
    port map (
            O => \N__33251\,
            I => \current_shift_inst.control_input_cry_28\
        );

    \I__6295\ : InMux
    port map (
            O => \N__33248\,
            I => \current_shift_inst.control_input_cry_29\
        );

    \I__6294\ : InMux
    port map (
            O => \N__33245\,
            I => \N__33242\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__33242\,
            I => \N__33238\
        );

    \I__6292\ : InMux
    port map (
            O => \N__33241\,
            I => \N__33235\
        );

    \I__6291\ : Odrv4
    port map (
            O => \N__33238\,
            I => \current_shift_inst.control_input_31\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__33235\,
            I => \current_shift_inst.control_input_31\
        );

    \I__6289\ : InMux
    port map (
            O => \N__33230\,
            I => \N__33227\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__33227\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\
        );

    \I__6287\ : IoInMux
    port map (
            O => \N__33224\,
            I => \N__33221\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__33221\,
            I => \N__33218\
        );

    \I__6285\ : Span4Mux_s0_v
    port map (
            O => \N__33218\,
            I => \N__33215\
        );

    \I__6284\ : Odrv4
    port map (
            O => \N__33215\,
            I => \pll_inst.red_c_i\
        );

    \I__6283\ : InMux
    port map (
            O => \N__33212\,
            I => \N__33208\
        );

    \I__6282\ : InMux
    port map (
            O => \N__33211\,
            I => \N__33204\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__33208\,
            I => \N__33201\
        );

    \I__6280\ : InMux
    port map (
            O => \N__33207\,
            I => \N__33198\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__33204\,
            I => \N__33195\
        );

    \I__6278\ : Span4Mux_v
    port map (
            O => \N__33201\,
            I => \N__33190\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__33198\,
            I => \N__33190\
        );

    \I__6276\ : Span12Mux_h
    port map (
            O => \N__33195\,
            I => \N__33187\
        );

    \I__6275\ : Span4Mux_h
    port map (
            O => \N__33190\,
            I => \N__33184\
        );

    \I__6274\ : Span12Mux_v
    port map (
            O => \N__33187\,
            I => \N__33181\
        );

    \I__6273\ : Span4Mux_v
    port map (
            O => \N__33184\,
            I => \N__33178\
        );

    \I__6272\ : Odrv12
    port map (
            O => \N__33181\,
            I => il_min_comp1_c
        );

    \I__6271\ : Odrv4
    port map (
            O => \N__33178\,
            I => il_min_comp1_c
        );

    \I__6270\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33170\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__33170\,
            I => \N__33167\
        );

    \I__6268\ : Odrv4
    port map (
            O => \N__33167\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\
        );

    \I__6267\ : InMux
    port map (
            O => \N__33164\,
            I => \current_shift_inst.control_input_cry_16\
        );

    \I__6266\ : CascadeMux
    port map (
            O => \N__33161\,
            I => \N__33158\
        );

    \I__6265\ : InMux
    port map (
            O => \N__33158\,
            I => \N__33155\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__33155\,
            I => \N__33152\
        );

    \I__6263\ : Odrv4
    port map (
            O => \N__33152\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\
        );

    \I__6262\ : InMux
    port map (
            O => \N__33149\,
            I => \current_shift_inst.control_input_cry_17\
        );

    \I__6261\ : InMux
    port map (
            O => \N__33146\,
            I => \N__33143\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__33143\,
            I => \N__33140\
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__33140\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\
        );

    \I__6258\ : InMux
    port map (
            O => \N__33137\,
            I => \current_shift_inst.control_input_cry_18\
        );

    \I__6257\ : InMux
    port map (
            O => \N__33134\,
            I => \N__33131\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__33131\,
            I => \N__33128\
        );

    \I__6255\ : Odrv4
    port map (
            O => \N__33128\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\
        );

    \I__6254\ : InMux
    port map (
            O => \N__33125\,
            I => \current_shift_inst.control_input_cry_19\
        );

    \I__6253\ : CascadeMux
    port map (
            O => \N__33122\,
            I => \N__33119\
        );

    \I__6252\ : InMux
    port map (
            O => \N__33119\,
            I => \N__33116\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__33116\,
            I => \N__33113\
        );

    \I__6250\ : Odrv4
    port map (
            O => \N__33113\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\
        );

    \I__6249\ : InMux
    port map (
            O => \N__33110\,
            I => \current_shift_inst.control_input_cry_20\
        );

    \I__6248\ : InMux
    port map (
            O => \N__33107\,
            I => \N__33104\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__33104\,
            I => \N__33101\
        );

    \I__6246\ : Odrv4
    port map (
            O => \N__33101\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\
        );

    \I__6245\ : InMux
    port map (
            O => \N__33098\,
            I => \current_shift_inst.control_input_cry_21\
        );

    \I__6244\ : CascadeMux
    port map (
            O => \N__33095\,
            I => \N__33092\
        );

    \I__6243\ : InMux
    port map (
            O => \N__33092\,
            I => \N__33089\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__33089\,
            I => \N__33086\
        );

    \I__6241\ : Odrv4
    port map (
            O => \N__33086\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\
        );

    \I__6240\ : InMux
    port map (
            O => \N__33083\,
            I => \current_shift_inst.control_input_cry_22\
        );

    \I__6239\ : CascadeMux
    port map (
            O => \N__33080\,
            I => \N__33077\
        );

    \I__6238\ : InMux
    port map (
            O => \N__33077\,
            I => \N__33074\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__33074\,
            I => \N__33071\
        );

    \I__6236\ : Odrv4
    port map (
            O => \N__33071\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\
        );

    \I__6235\ : InMux
    port map (
            O => \N__33068\,
            I => \bfn_12_20_0_\
        );

    \I__6234\ : CascadeMux
    port map (
            O => \N__33065\,
            I => \N__33062\
        );

    \I__6233\ : InMux
    port map (
            O => \N__33062\,
            I => \N__33059\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__33059\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__6231\ : InMux
    port map (
            O => \N__33056\,
            I => \N__33053\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__33053\,
            I => \N__33050\
        );

    \I__6229\ : Odrv4
    port map (
            O => \N__33050\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__6228\ : InMux
    port map (
            O => \N__33047\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__6227\ : CascadeMux
    port map (
            O => \N__33044\,
            I => \N__33041\
        );

    \I__6226\ : InMux
    port map (
            O => \N__33041\,
            I => \N__33038\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__33038\,
            I => \N__33035\
        );

    \I__6224\ : Odrv4
    port map (
            O => \N__33035\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__6223\ : InMux
    port map (
            O => \N__33032\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__6222\ : InMux
    port map (
            O => \N__33029\,
            I => \N__33026\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__33026\,
            I => \N__33023\
        );

    \I__6220\ : Odrv4
    port map (
            O => \N__33023\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__6219\ : InMux
    port map (
            O => \N__33020\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__6218\ : InMux
    port map (
            O => \N__33017\,
            I => \N__33014\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__33014\,
            I => \N__33011\
        );

    \I__6216\ : Odrv4
    port map (
            O => \N__33011\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__6215\ : InMux
    port map (
            O => \N__33008\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__6214\ : CascadeMux
    port map (
            O => \N__33005\,
            I => \N__33002\
        );

    \I__6213\ : InMux
    port map (
            O => \N__33002\,
            I => \N__32999\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__32999\,
            I => \N__32996\
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__32996\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__6210\ : InMux
    port map (
            O => \N__32993\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__6209\ : InMux
    port map (
            O => \N__32990\,
            I => \N__32987\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__32987\,
            I => \N__32984\
        );

    \I__6207\ : Odrv4
    port map (
            O => \N__32984\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\
        );

    \I__6206\ : InMux
    port map (
            O => \N__32981\,
            I => \current_shift_inst.control_input_cry_13\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__32978\,
            I => \N__32975\
        );

    \I__6204\ : InMux
    port map (
            O => \N__32975\,
            I => \N__32972\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__32972\,
            I => \N__32969\
        );

    \I__6202\ : Odrv4
    port map (
            O => \N__32969\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\
        );

    \I__6201\ : InMux
    port map (
            O => \N__32966\,
            I => \current_shift_inst.control_input_cry_14\
        );

    \I__6200\ : CascadeMux
    port map (
            O => \N__32963\,
            I => \N__32960\
        );

    \I__6199\ : InMux
    port map (
            O => \N__32960\,
            I => \N__32957\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__32957\,
            I => \N__32954\
        );

    \I__6197\ : Odrv4
    port map (
            O => \N__32954\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\
        );

    \I__6196\ : InMux
    port map (
            O => \N__32951\,
            I => \bfn_12_19_0_\
        );

    \I__6195\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32945\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__32945\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__6193\ : CascadeMux
    port map (
            O => \N__32942\,
            I => \N__32939\
        );

    \I__6192\ : InMux
    port map (
            O => \N__32939\,
            I => \N__32936\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__32936\,
            I => \N__32931\
        );

    \I__6190\ : InMux
    port map (
            O => \N__32935\,
            I => \N__32928\
        );

    \I__6189\ : InMux
    port map (
            O => \N__32934\,
            I => \N__32925\
        );

    \I__6188\ : Span4Mux_h
    port map (
            O => \N__32931\,
            I => \N__32922\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__32928\,
            I => \current_shift_inst.N_1271_i\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__32925\,
            I => \current_shift_inst.N_1271_i\
        );

    \I__6185\ : Odrv4
    port map (
            O => \N__32922\,
            I => \current_shift_inst.N_1271_i\
        );

    \I__6184\ : InMux
    port map (
            O => \N__32915\,
            I => \N__32912\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__32912\,
            I => \N__32909\
        );

    \I__6182\ : Odrv4
    port map (
            O => \N__32909\,
            I => \current_shift_inst.control_input_1\
        );

    \I__6181\ : InMux
    port map (
            O => \N__32906\,
            I => \N__32903\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__32903\,
            I => \N__32900\
        );

    \I__6179\ : Odrv4
    port map (
            O => \N__32900\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__6178\ : InMux
    port map (
            O => \N__32897\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__6177\ : CascadeMux
    port map (
            O => \N__32894\,
            I => \N__32891\
        );

    \I__6176\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32888\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__32888\,
            I => \N__32885\
        );

    \I__6174\ : Odrv4
    port map (
            O => \N__32885\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__6173\ : InMux
    port map (
            O => \N__32882\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__6172\ : InMux
    port map (
            O => \N__32879\,
            I => \N__32876\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__32876\,
            I => \N__32873\
        );

    \I__6170\ : Odrv4
    port map (
            O => \N__32873\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__6169\ : InMux
    port map (
            O => \N__32870\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__6168\ : InMux
    port map (
            O => \N__32867\,
            I => \N__32864\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__32864\,
            I => \N__32861\
        );

    \I__6166\ : Odrv4
    port map (
            O => \N__32861\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__6165\ : InMux
    port map (
            O => \N__32858\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__6164\ : CascadeMux
    port map (
            O => \N__32855\,
            I => \N__32852\
        );

    \I__6163\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32849\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__32849\,
            I => \N__32846\
        );

    \I__6161\ : Odrv4
    port map (
            O => \N__32846\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__6160\ : InMux
    port map (
            O => \N__32843\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__6159\ : InMux
    port map (
            O => \N__32840\,
            I => \N__32837\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__32837\,
            I => \N__32834\
        );

    \I__6157\ : Odrv4
    port map (
            O => \N__32834\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__6156\ : InMux
    port map (
            O => \N__32831\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__6155\ : CascadeMux
    port map (
            O => \N__32828\,
            I => \N__32825\
        );

    \I__6154\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32822\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__32822\,
            I => \N__32819\
        );

    \I__6152\ : Odrv4
    port map (
            O => \N__32819\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__6151\ : InMux
    port map (
            O => \N__32816\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__6150\ : InMux
    port map (
            O => \N__32813\,
            I => \N__32810\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__32810\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__6148\ : CascadeMux
    port map (
            O => \N__32807\,
            I => \N__32804\
        );

    \I__6147\ : InMux
    port map (
            O => \N__32804\,
            I => \N__32801\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__32801\,
            I => \N__32798\
        );

    \I__6145\ : Odrv4
    port map (
            O => \N__32798\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__6144\ : InMux
    port map (
            O => \N__32795\,
            I => \bfn_12_18_0_\
        );

    \I__6143\ : InMux
    port map (
            O => \N__32792\,
            I => \N__32785\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32791\,
            I => \N__32785\
        );

    \I__6141\ : InMux
    port map (
            O => \N__32790\,
            I => \N__32782\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__32785\,
            I => \N__32779\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__32782\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__6138\ : Odrv4
    port map (
            O => \N__32779\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__6137\ : InMux
    port map (
            O => \N__32774\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__6136\ : CascadeMux
    port map (
            O => \N__32771\,
            I => \N__32767\
        );

    \I__6135\ : CascadeMux
    port map (
            O => \N__32770\,
            I => \N__32764\
        );

    \I__6134\ : InMux
    port map (
            O => \N__32767\,
            I => \N__32761\
        );

    \I__6133\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32757\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__32761\,
            I => \N__32754\
        );

    \I__6131\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32751\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__32757\,
            I => \N__32746\
        );

    \I__6129\ : Span4Mux_h
    port map (
            O => \N__32754\,
            I => \N__32746\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__32751\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__6127\ : Odrv4
    port map (
            O => \N__32746\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__6126\ : InMux
    port map (
            O => \N__32741\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__6125\ : CEMux
    port map (
            O => \N__32738\,
            I => \N__32733\
        );

    \I__6124\ : CEMux
    port map (
            O => \N__32737\,
            I => \N__32730\
        );

    \I__6123\ : CEMux
    port map (
            O => \N__32736\,
            I => \N__32727\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__32733\,
            I => \N__32716\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__32730\,
            I => \N__32716\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__32727\,
            I => \N__32699\
        );

    \I__6119\ : CEMux
    port map (
            O => \N__32726\,
            I => \N__32696\
        );

    \I__6118\ : CEMux
    port map (
            O => \N__32725\,
            I => \N__32693\
        );

    \I__6117\ : InMux
    port map (
            O => \N__32724\,
            I => \N__32680\
        );

    \I__6116\ : InMux
    port map (
            O => \N__32723\,
            I => \N__32680\
        );

    \I__6115\ : InMux
    port map (
            O => \N__32722\,
            I => \N__32680\
        );

    \I__6114\ : CEMux
    port map (
            O => \N__32721\,
            I => \N__32676\
        );

    \I__6113\ : Span4Mux_v
    port map (
            O => \N__32716\,
            I => \N__32662\
        );

    \I__6112\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32653\
        );

    \I__6111\ : InMux
    port map (
            O => \N__32714\,
            I => \N__32653\
        );

    \I__6110\ : InMux
    port map (
            O => \N__32713\,
            I => \N__32653\
        );

    \I__6109\ : InMux
    port map (
            O => \N__32712\,
            I => \N__32653\
        );

    \I__6108\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32644\
        );

    \I__6107\ : InMux
    port map (
            O => \N__32710\,
            I => \N__32644\
        );

    \I__6106\ : InMux
    port map (
            O => \N__32709\,
            I => \N__32644\
        );

    \I__6105\ : InMux
    port map (
            O => \N__32708\,
            I => \N__32644\
        );

    \I__6104\ : InMux
    port map (
            O => \N__32707\,
            I => \N__32635\
        );

    \I__6103\ : InMux
    port map (
            O => \N__32706\,
            I => \N__32635\
        );

    \I__6102\ : InMux
    port map (
            O => \N__32705\,
            I => \N__32635\
        );

    \I__6101\ : InMux
    port map (
            O => \N__32704\,
            I => \N__32635\
        );

    \I__6100\ : CEMux
    port map (
            O => \N__32703\,
            I => \N__32632\
        );

    \I__6099\ : CEMux
    port map (
            O => \N__32702\,
            I => \N__32628\
        );

    \I__6098\ : Span4Mux_v
    port map (
            O => \N__32699\,
            I => \N__32620\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__32696\,
            I => \N__32620\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__32693\,
            I => \N__32620\
        );

    \I__6095\ : InMux
    port map (
            O => \N__32692\,
            I => \N__32611\
        );

    \I__6094\ : InMux
    port map (
            O => \N__32691\,
            I => \N__32611\
        );

    \I__6093\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32611\
        );

    \I__6092\ : InMux
    port map (
            O => \N__32689\,
            I => \N__32611\
        );

    \I__6091\ : InMux
    port map (
            O => \N__32688\,
            I => \N__32608\
        );

    \I__6090\ : CEMux
    port map (
            O => \N__32687\,
            I => \N__32605\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__32680\,
            I => \N__32602\
        );

    \I__6088\ : CEMux
    port map (
            O => \N__32679\,
            I => \N__32599\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__32676\,
            I => \N__32596\
        );

    \I__6086\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32587\
        );

    \I__6085\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32587\
        );

    \I__6084\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32587\
        );

    \I__6083\ : InMux
    port map (
            O => \N__32672\,
            I => \N__32587\
        );

    \I__6082\ : InMux
    port map (
            O => \N__32671\,
            I => \N__32580\
        );

    \I__6081\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32580\
        );

    \I__6080\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32580\
        );

    \I__6079\ : InMux
    port map (
            O => \N__32668\,
            I => \N__32571\
        );

    \I__6078\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32571\
        );

    \I__6077\ : InMux
    port map (
            O => \N__32666\,
            I => \N__32571\
        );

    \I__6076\ : InMux
    port map (
            O => \N__32665\,
            I => \N__32571\
        );

    \I__6075\ : Span4Mux_v
    port map (
            O => \N__32662\,
            I => \N__32564\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__32653\,
            I => \N__32564\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__32644\,
            I => \N__32564\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__32635\,
            I => \N__32561\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__32632\,
            I => \N__32557\
        );

    \I__6070\ : CEMux
    port map (
            O => \N__32631\,
            I => \N__32554\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__32628\,
            I => \N__32551\
        );

    \I__6068\ : CEMux
    port map (
            O => \N__32627\,
            I => \N__32548\
        );

    \I__6067\ : Span4Mux_h
    port map (
            O => \N__32620\,
            I => \N__32545\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__32611\,
            I => \N__32542\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__32608\,
            I => \N__32539\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__32605\,
            I => \N__32534\
        );

    \I__6063\ : Span4Mux_h
    port map (
            O => \N__32602\,
            I => \N__32534\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__32599\,
            I => \N__32529\
        );

    \I__6061\ : Span4Mux_v
    port map (
            O => \N__32596\,
            I => \N__32529\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__32587\,
            I => \N__32518\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__32580\,
            I => \N__32518\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__32571\,
            I => \N__32518\
        );

    \I__6057\ : Span4Mux_h
    port map (
            O => \N__32564\,
            I => \N__32518\
        );

    \I__6056\ : Span4Mux_v
    port map (
            O => \N__32561\,
            I => \N__32518\
        );

    \I__6055\ : CEMux
    port map (
            O => \N__32560\,
            I => \N__32515\
        );

    \I__6054\ : Span4Mux_v
    port map (
            O => \N__32557\,
            I => \N__32512\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__32554\,
            I => \N__32507\
        );

    \I__6052\ : Sp12to4
    port map (
            O => \N__32551\,
            I => \N__32507\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__32548\,
            I => \N__32500\
        );

    \I__6050\ : Span4Mux_v
    port map (
            O => \N__32545\,
            I => \N__32500\
        );

    \I__6049\ : Span4Mux_h
    port map (
            O => \N__32542\,
            I => \N__32500\
        );

    \I__6048\ : Span4Mux_h
    port map (
            O => \N__32539\,
            I => \N__32495\
        );

    \I__6047\ : Span4Mux_v
    port map (
            O => \N__32534\,
            I => \N__32495\
        );

    \I__6046\ : Span4Mux_v
    port map (
            O => \N__32529\,
            I => \N__32490\
        );

    \I__6045\ : Span4Mux_v
    port map (
            O => \N__32518\,
            I => \N__32490\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__32515\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__32512\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6042\ : Odrv12
    port map (
            O => \N__32507\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6041\ : Odrv4
    port map (
            O => \N__32500\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__32495\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6039\ : Odrv4
    port map (
            O => \N__32490\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6038\ : InMux
    port map (
            O => \N__32477\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__6037\ : InMux
    port map (
            O => \N__32474\,
            I => \N__32469\
        );

    \I__6036\ : InMux
    port map (
            O => \N__32473\,
            I => \N__32466\
        );

    \I__6035\ : InMux
    port map (
            O => \N__32472\,
            I => \N__32463\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__32469\,
            I => \N__32458\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__32466\,
            I => \N__32458\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__32463\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__6031\ : Odrv12
    port map (
            O => \N__32458\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__6030\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32450\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__32450\,
            I => \N__32445\
        );

    \I__6028\ : InMux
    port map (
            O => \N__32449\,
            I => \N__32442\
        );

    \I__6027\ : InMux
    port map (
            O => \N__32448\,
            I => \N__32439\
        );

    \I__6026\ : Span4Mux_h
    port map (
            O => \N__32445\,
            I => \N__32436\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__32442\,
            I => \N__32433\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__32439\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__6023\ : Odrv4
    port map (
            O => \N__32436\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__6022\ : Odrv12
    port map (
            O => \N__32433\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__6021\ : InMux
    port map (
            O => \N__32426\,
            I => \N__32387\
        );

    \I__6020\ : InMux
    port map (
            O => \N__32425\,
            I => \N__32387\
        );

    \I__6019\ : InMux
    port map (
            O => \N__32424\,
            I => \N__32380\
        );

    \I__6018\ : InMux
    port map (
            O => \N__32423\,
            I => \N__32380\
        );

    \I__6017\ : InMux
    port map (
            O => \N__32422\,
            I => \N__32380\
        );

    \I__6016\ : InMux
    port map (
            O => \N__32421\,
            I => \N__32373\
        );

    \I__6015\ : InMux
    port map (
            O => \N__32420\,
            I => \N__32373\
        );

    \I__6014\ : InMux
    port map (
            O => \N__32419\,
            I => \N__32373\
        );

    \I__6013\ : InMux
    port map (
            O => \N__32418\,
            I => \N__32368\
        );

    \I__6012\ : InMux
    port map (
            O => \N__32417\,
            I => \N__32368\
        );

    \I__6011\ : InMux
    port map (
            O => \N__32416\,
            I => \N__32363\
        );

    \I__6010\ : InMux
    port map (
            O => \N__32415\,
            I => \N__32363\
        );

    \I__6009\ : InMux
    port map (
            O => \N__32414\,
            I => \N__32341\
        );

    \I__6008\ : InMux
    port map (
            O => \N__32413\,
            I => \N__32319\
        );

    \I__6007\ : InMux
    port map (
            O => \N__32412\,
            I => \N__32319\
        );

    \I__6006\ : InMux
    port map (
            O => \N__32411\,
            I => \N__32316\
        );

    \I__6005\ : InMux
    port map (
            O => \N__32410\,
            I => \N__32313\
        );

    \I__6004\ : InMux
    port map (
            O => \N__32409\,
            I => \N__32310\
        );

    \I__6003\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32300\
        );

    \I__6002\ : InMux
    port map (
            O => \N__32407\,
            I => \N__32291\
        );

    \I__6001\ : InMux
    port map (
            O => \N__32406\,
            I => \N__32291\
        );

    \I__6000\ : InMux
    port map (
            O => \N__32405\,
            I => \N__32291\
        );

    \I__5999\ : InMux
    port map (
            O => \N__32404\,
            I => \N__32291\
        );

    \I__5998\ : InMux
    port map (
            O => \N__32403\,
            I => \N__32278\
        );

    \I__5997\ : InMux
    port map (
            O => \N__32402\,
            I => \N__32278\
        );

    \I__5996\ : InMux
    port map (
            O => \N__32401\,
            I => \N__32278\
        );

    \I__5995\ : InMux
    port map (
            O => \N__32400\,
            I => \N__32278\
        );

    \I__5994\ : InMux
    port map (
            O => \N__32399\,
            I => \N__32278\
        );

    \I__5993\ : InMux
    port map (
            O => \N__32398\,
            I => \N__32278\
        );

    \I__5992\ : InMux
    port map (
            O => \N__32397\,
            I => \N__32269\
        );

    \I__5991\ : InMux
    port map (
            O => \N__32396\,
            I => \N__32269\
        );

    \I__5990\ : InMux
    port map (
            O => \N__32395\,
            I => \N__32269\
        );

    \I__5989\ : InMux
    port map (
            O => \N__32394\,
            I => \N__32269\
        );

    \I__5988\ : InMux
    port map (
            O => \N__32393\,
            I => \N__32264\
        );

    \I__5987\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32264\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__32387\,
            I => \N__32253\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__32380\,
            I => \N__32253\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__32373\,
            I => \N__32253\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__32368\,
            I => \N__32253\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__32363\,
            I => \N__32253\
        );

    \I__5981\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32242\
        );

    \I__5980\ : InMux
    port map (
            O => \N__32361\,
            I => \N__32242\
        );

    \I__5979\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32242\
        );

    \I__5978\ : InMux
    port map (
            O => \N__32359\,
            I => \N__32242\
        );

    \I__5977\ : InMux
    port map (
            O => \N__32358\,
            I => \N__32242\
        );

    \I__5976\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32239\
        );

    \I__5975\ : InMux
    port map (
            O => \N__32356\,
            I => \N__32228\
        );

    \I__5974\ : InMux
    port map (
            O => \N__32355\,
            I => \N__32228\
        );

    \I__5973\ : InMux
    port map (
            O => \N__32354\,
            I => \N__32228\
        );

    \I__5972\ : InMux
    port map (
            O => \N__32353\,
            I => \N__32228\
        );

    \I__5971\ : InMux
    port map (
            O => \N__32352\,
            I => \N__32228\
        );

    \I__5970\ : InMux
    port map (
            O => \N__32351\,
            I => \N__32217\
        );

    \I__5969\ : InMux
    port map (
            O => \N__32350\,
            I => \N__32217\
        );

    \I__5968\ : InMux
    port map (
            O => \N__32349\,
            I => \N__32217\
        );

    \I__5967\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32217\
        );

    \I__5966\ : InMux
    port map (
            O => \N__32347\,
            I => \N__32217\
        );

    \I__5965\ : InMux
    port map (
            O => \N__32346\,
            I => \N__32210\
        );

    \I__5964\ : InMux
    port map (
            O => \N__32345\,
            I => \N__32210\
        );

    \I__5963\ : InMux
    port map (
            O => \N__32344\,
            I => \N__32210\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__32341\,
            I => \N__32207\
        );

    \I__5961\ : InMux
    port map (
            O => \N__32340\,
            I => \N__32200\
        );

    \I__5960\ : InMux
    port map (
            O => \N__32339\,
            I => \N__32200\
        );

    \I__5959\ : InMux
    port map (
            O => \N__32338\,
            I => \N__32200\
        );

    \I__5958\ : InMux
    port map (
            O => \N__32337\,
            I => \N__32191\
        );

    \I__5957\ : InMux
    port map (
            O => \N__32336\,
            I => \N__32191\
        );

    \I__5956\ : InMux
    port map (
            O => \N__32335\,
            I => \N__32191\
        );

    \I__5955\ : InMux
    port map (
            O => \N__32334\,
            I => \N__32191\
        );

    \I__5954\ : InMux
    port map (
            O => \N__32333\,
            I => \N__32171\
        );

    \I__5953\ : InMux
    port map (
            O => \N__32332\,
            I => \N__32171\
        );

    \I__5952\ : InMux
    port map (
            O => \N__32331\,
            I => \N__32171\
        );

    \I__5951\ : InMux
    port map (
            O => \N__32330\,
            I => \N__32171\
        );

    \I__5950\ : InMux
    port map (
            O => \N__32329\,
            I => \N__32171\
        );

    \I__5949\ : InMux
    port map (
            O => \N__32328\,
            I => \N__32171\
        );

    \I__5948\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32161\
        );

    \I__5947\ : InMux
    port map (
            O => \N__32326\,
            I => \N__32156\
        );

    \I__5946\ : InMux
    port map (
            O => \N__32325\,
            I => \N__32156\
        );

    \I__5945\ : InMux
    port map (
            O => \N__32324\,
            I => \N__32153\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__32319\,
            I => \N__32150\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__32316\,
            I => \N__32143\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__32313\,
            I => \N__32143\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__32310\,
            I => \N__32143\
        );

    \I__5940\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32128\
        );

    \I__5939\ : InMux
    port map (
            O => \N__32308\,
            I => \N__32128\
        );

    \I__5938\ : InMux
    port map (
            O => \N__32307\,
            I => \N__32128\
        );

    \I__5937\ : InMux
    port map (
            O => \N__32306\,
            I => \N__32128\
        );

    \I__5936\ : InMux
    port map (
            O => \N__32305\,
            I => \N__32128\
        );

    \I__5935\ : InMux
    port map (
            O => \N__32304\,
            I => \N__32128\
        );

    \I__5934\ : InMux
    port map (
            O => \N__32303\,
            I => \N__32128\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__32300\,
            I => \N__32115\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__32291\,
            I => \N__32115\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__32278\,
            I => \N__32115\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__32269\,
            I => \N__32115\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__32264\,
            I => \N__32115\
        );

    \I__5928\ : Span4Mux_v
    port map (
            O => \N__32253\,
            I => \N__32115\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__32242\,
            I => \N__32112\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__32239\,
            I => \N__32107\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__32228\,
            I => \N__32107\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__32217\,
            I => \N__32096\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__32210\,
            I => \N__32096\
        );

    \I__5922\ : Span4Mux_v
    port map (
            O => \N__32207\,
            I => \N__32096\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__32200\,
            I => \N__32096\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__32191\,
            I => \N__32096\
        );

    \I__5919\ : InMux
    port map (
            O => \N__32190\,
            I => \N__32093\
        );

    \I__5918\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32090\
        );

    \I__5917\ : InMux
    port map (
            O => \N__32188\,
            I => \N__32079\
        );

    \I__5916\ : InMux
    port map (
            O => \N__32187\,
            I => \N__32079\
        );

    \I__5915\ : InMux
    port map (
            O => \N__32186\,
            I => \N__32079\
        );

    \I__5914\ : InMux
    port map (
            O => \N__32185\,
            I => \N__32079\
        );

    \I__5913\ : InMux
    port map (
            O => \N__32184\,
            I => \N__32079\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__32171\,
            I => \N__32076\
        );

    \I__5911\ : InMux
    port map (
            O => \N__32170\,
            I => \N__32067\
        );

    \I__5910\ : InMux
    port map (
            O => \N__32169\,
            I => \N__32067\
        );

    \I__5909\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32067\
        );

    \I__5908\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32067\
        );

    \I__5907\ : InMux
    port map (
            O => \N__32166\,
            I => \N__32062\
        );

    \I__5906\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32062\
        );

    \I__5905\ : InMux
    port map (
            O => \N__32164\,
            I => \N__32059\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__32161\,
            I => \N__32054\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__32156\,
            I => \N__32054\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__32153\,
            I => \N__32051\
        );

    \I__5901\ : Span4Mux_v
    port map (
            O => \N__32150\,
            I => \N__32048\
        );

    \I__5900\ : Span4Mux_v
    port map (
            O => \N__32143\,
            I => \N__32041\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__32128\,
            I => \N__32041\
        );

    \I__5898\ : Span4Mux_v
    port map (
            O => \N__32115\,
            I => \N__32041\
        );

    \I__5897\ : Span12Mux_s11_h
    port map (
            O => \N__32112\,
            I => \N__32038\
        );

    \I__5896\ : Span4Mux_h
    port map (
            O => \N__32107\,
            I => \N__32033\
        );

    \I__5895\ : Span4Mux_v
    port map (
            O => \N__32096\,
            I => \N__32033\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__32093\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__32090\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__32079\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__32076\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__32067\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__32062\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__32059\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5887\ : Odrv4
    port map (
            O => \N__32054\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5886\ : Odrv4
    port map (
            O => \N__32051\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5885\ : Odrv4
    port map (
            O => \N__32048\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5884\ : Odrv4
    port map (
            O => \N__32041\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5883\ : Odrv12
    port map (
            O => \N__32038\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5882\ : Odrv4
    port map (
            O => \N__32033\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5881\ : InMux
    port map (
            O => \N__32006\,
            I => \N__32003\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__32003\,
            I => \N__31998\
        );

    \I__5879\ : InMux
    port map (
            O => \N__32002\,
            I => \N__31995\
        );

    \I__5878\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31992\
        );

    \I__5877\ : Span4Mux_h
    port map (
            O => \N__31998\,
            I => \N__31989\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__31995\,
            I => \N__31986\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__31992\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__5874\ : Odrv4
    port map (
            O => \N__31989\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__5873\ : Odrv4
    port map (
            O => \N__31986\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__5872\ : InMux
    port map (
            O => \N__31979\,
            I => \N__31976\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__31976\,
            I => \N__31972\
        );

    \I__5870\ : InMux
    port map (
            O => \N__31975\,
            I => \N__31969\
        );

    \I__5869\ : Odrv12
    port map (
            O => \N__31972\,
            I => \phase_controller_inst1.N_52\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__31969\,
            I => \phase_controller_inst1.N_52\
        );

    \I__5867\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31961\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__31961\,
            I => \phase_controller_inst1_N_54\
        );

    \I__5865\ : CascadeMux
    port map (
            O => \N__31958\,
            I => \N__31955\
        );

    \I__5864\ : InMux
    port map (
            O => \N__31955\,
            I => \N__31951\
        );

    \I__5863\ : InMux
    port map (
            O => \N__31954\,
            I => \N__31947\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__31951\,
            I => \N__31942\
        );

    \I__5861\ : InMux
    port map (
            O => \N__31950\,
            I => \N__31939\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__31947\,
            I => \N__31936\
        );

    \I__5859\ : InMux
    port map (
            O => \N__31946\,
            I => \N__31933\
        );

    \I__5858\ : InMux
    port map (
            O => \N__31945\,
            I => \N__31930\
        );

    \I__5857\ : Span4Mux_v
    port map (
            O => \N__31942\,
            I => \N__31925\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__31939\,
            I => \N__31925\
        );

    \I__5855\ : Span4Mux_v
    port map (
            O => \N__31936\,
            I => \N__31922\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__31933\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__31930\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__5852\ : Odrv4
    port map (
            O => \N__31925\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__5851\ : Odrv4
    port map (
            O => \N__31922\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__5850\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31909\
        );

    \I__5849\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31906\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__31909\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__31906\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__5846\ : InMux
    port map (
            O => \N__31901\,
            I => \N__31897\
        );

    \I__5845\ : InMux
    port map (
            O => \N__31900\,
            I => \N__31893\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__31897\,
            I => \N__31890\
        );

    \I__5843\ : InMux
    port map (
            O => \N__31896\,
            I => \N__31887\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__31893\,
            I => \N__31884\
        );

    \I__5841\ : Span4Mux_h
    port map (
            O => \N__31890\,
            I => \N__31881\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__31887\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__5839\ : Odrv4
    port map (
            O => \N__31884\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__5838\ : Odrv4
    port map (
            O => \N__31881\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__5837\ : InMux
    port map (
            O => \N__31874\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__5836\ : InMux
    port map (
            O => \N__31871\,
            I => \N__31867\
        );

    \I__5835\ : InMux
    port map (
            O => \N__31870\,
            I => \N__31863\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__31867\,
            I => \N__31860\
        );

    \I__5833\ : InMux
    port map (
            O => \N__31866\,
            I => \N__31857\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__31863\,
            I => \N__31852\
        );

    \I__5831\ : Span4Mux_v
    port map (
            O => \N__31860\,
            I => \N__31852\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__31857\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__5829\ : Odrv4
    port map (
            O => \N__31852\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__5828\ : InMux
    port map (
            O => \N__31847\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__5827\ : InMux
    port map (
            O => \N__31844\,
            I => \N__31838\
        );

    \I__5826\ : InMux
    port map (
            O => \N__31843\,
            I => \N__31838\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__31838\,
            I => \N__31834\
        );

    \I__5824\ : InMux
    port map (
            O => \N__31837\,
            I => \N__31831\
        );

    \I__5823\ : Span4Mux_h
    port map (
            O => \N__31834\,
            I => \N__31828\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__31831\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__31828\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__5820\ : InMux
    port map (
            O => \N__31823\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__5819\ : CascadeMux
    port map (
            O => \N__31820\,
            I => \N__31816\
        );

    \I__5818\ : CascadeMux
    port map (
            O => \N__31819\,
            I => \N__31813\
        );

    \I__5817\ : InMux
    port map (
            O => \N__31816\,
            I => \N__31810\
        );

    \I__5816\ : InMux
    port map (
            O => \N__31813\,
            I => \N__31807\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__31810\,
            I => \N__31801\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__31807\,
            I => \N__31801\
        );

    \I__5813\ : InMux
    port map (
            O => \N__31806\,
            I => \N__31798\
        );

    \I__5812\ : Span12Mux_s11_v
    port map (
            O => \N__31801\,
            I => \N__31795\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__31798\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__5810\ : Odrv12
    port map (
            O => \N__31795\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__5809\ : InMux
    port map (
            O => \N__31790\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__5808\ : CascadeMux
    port map (
            O => \N__31787\,
            I => \N__31783\
        );

    \I__5807\ : CascadeMux
    port map (
            O => \N__31786\,
            I => \N__31780\
        );

    \I__5806\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31774\
        );

    \I__5805\ : InMux
    port map (
            O => \N__31780\,
            I => \N__31774\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31779\,
            I => \N__31771\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__31774\,
            I => \N__31768\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__31771\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__5801\ : Odrv4
    port map (
            O => \N__31768\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__5800\ : InMux
    port map (
            O => \N__31763\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__5799\ : InMux
    port map (
            O => \N__31760\,
            I => \N__31754\
        );

    \I__5798\ : InMux
    port map (
            O => \N__31759\,
            I => \N__31754\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__31754\,
            I => \N__31750\
        );

    \I__5796\ : InMux
    port map (
            O => \N__31753\,
            I => \N__31747\
        );

    \I__5795\ : Span4Mux_v
    port map (
            O => \N__31750\,
            I => \N__31744\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__31747\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__5793\ : Odrv4
    port map (
            O => \N__31744\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__5792\ : InMux
    port map (
            O => \N__31739\,
            I => \bfn_12_13_0_\
        );

    \I__5791\ : CascadeMux
    port map (
            O => \N__31736\,
            I => \N__31733\
        );

    \I__5790\ : InMux
    port map (
            O => \N__31733\,
            I => \N__31726\
        );

    \I__5789\ : InMux
    port map (
            O => \N__31732\,
            I => \N__31726\
        );

    \I__5788\ : InMux
    port map (
            O => \N__31731\,
            I => \N__31723\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__31726\,
            I => \N__31720\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__31723\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__5785\ : Odrv12
    port map (
            O => \N__31720\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__5784\ : InMux
    port map (
            O => \N__31715\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__5783\ : InMux
    port map (
            O => \N__31712\,
            I => \N__31705\
        );

    \I__5782\ : InMux
    port map (
            O => \N__31711\,
            I => \N__31705\
        );

    \I__5781\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31702\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__31705\,
            I => \N__31699\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__31702\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__5778\ : Odrv4
    port map (
            O => \N__31699\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__5777\ : InMux
    port map (
            O => \N__31694\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__5776\ : CascadeMux
    port map (
            O => \N__31691\,
            I => \N__31688\
        );

    \I__5775\ : InMux
    port map (
            O => \N__31688\,
            I => \N__31681\
        );

    \I__5774\ : InMux
    port map (
            O => \N__31687\,
            I => \N__31681\
        );

    \I__5773\ : InMux
    port map (
            O => \N__31686\,
            I => \N__31678\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__31681\,
            I => \N__31675\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__31678\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__5770\ : Odrv4
    port map (
            O => \N__31675\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__5769\ : InMux
    port map (
            O => \N__31670\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__5768\ : InMux
    port map (
            O => \N__31667\,
            I => \N__31664\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__31664\,
            I => \N__31660\
        );

    \I__5766\ : InMux
    port map (
            O => \N__31663\,
            I => \N__31657\
        );

    \I__5765\ : Span4Mux_h
    port map (
            O => \N__31660\,
            I => \N__31654\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__31657\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__5763\ : Odrv4
    port map (
            O => \N__31654\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__5762\ : InMux
    port map (
            O => \N__31649\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__5761\ : InMux
    port map (
            O => \N__31646\,
            I => \N__31643\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__31643\,
            I => \N__31639\
        );

    \I__5759\ : InMux
    port map (
            O => \N__31642\,
            I => \N__31636\
        );

    \I__5758\ : Span4Mux_h
    port map (
            O => \N__31639\,
            I => \N__31633\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__31636\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__5756\ : Odrv4
    port map (
            O => \N__31633\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__5755\ : InMux
    port map (
            O => \N__31628\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__5754\ : InMux
    port map (
            O => \N__31625\,
            I => \N__31622\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__31622\,
            I => \N__31618\
        );

    \I__5752\ : InMux
    port map (
            O => \N__31621\,
            I => \N__31615\
        );

    \I__5751\ : Span4Mux_h
    port map (
            O => \N__31618\,
            I => \N__31612\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__31615\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__5749\ : Odrv4
    port map (
            O => \N__31612\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__5748\ : InMux
    port map (
            O => \N__31607\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__5747\ : InMux
    port map (
            O => \N__31604\,
            I => \N__31601\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__31601\,
            I => \N__31597\
        );

    \I__5745\ : InMux
    port map (
            O => \N__31600\,
            I => \N__31594\
        );

    \I__5744\ : Span4Mux_h
    port map (
            O => \N__31597\,
            I => \N__31591\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__31594\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__5742\ : Odrv4
    port map (
            O => \N__31591\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__5741\ : InMux
    port map (
            O => \N__31586\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__5740\ : CascadeMux
    port map (
            O => \N__31583\,
            I => \N__31580\
        );

    \I__5739\ : InMux
    port map (
            O => \N__31580\,
            I => \N__31574\
        );

    \I__5738\ : InMux
    port map (
            O => \N__31579\,
            I => \N__31574\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__31574\,
            I => \N__31570\
        );

    \I__5736\ : InMux
    port map (
            O => \N__31573\,
            I => \N__31567\
        );

    \I__5735\ : Span4Mux_v
    port map (
            O => \N__31570\,
            I => \N__31564\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__31567\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__5733\ : Odrv4
    port map (
            O => \N__31564\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__5732\ : InMux
    port map (
            O => \N__31559\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__5731\ : InMux
    port map (
            O => \N__31556\,
            I => \N__31549\
        );

    \I__5730\ : InMux
    port map (
            O => \N__31555\,
            I => \N__31549\
        );

    \I__5729\ : InMux
    port map (
            O => \N__31554\,
            I => \N__31546\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__31549\,
            I => \N__31543\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__31546\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__5726\ : Odrv4
    port map (
            O => \N__31543\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__5725\ : InMux
    port map (
            O => \N__31538\,
            I => \bfn_12_12_0_\
        );

    \I__5724\ : InMux
    port map (
            O => \N__31535\,
            I => \N__31529\
        );

    \I__5723\ : InMux
    port map (
            O => \N__31534\,
            I => \N__31529\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__31529\,
            I => \N__31526\
        );

    \I__5721\ : Span4Mux_h
    port map (
            O => \N__31526\,
            I => \N__31522\
        );

    \I__5720\ : InMux
    port map (
            O => \N__31525\,
            I => \N__31519\
        );

    \I__5719\ : Span4Mux_v
    port map (
            O => \N__31522\,
            I => \N__31516\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__31519\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__5717\ : Odrv4
    port map (
            O => \N__31516\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__5716\ : InMux
    port map (
            O => \N__31511\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__5715\ : CascadeMux
    port map (
            O => \N__31508\,
            I => \N__31504\
        );

    \I__5714\ : InMux
    port map (
            O => \N__31507\,
            I => \N__31499\
        );

    \I__5713\ : InMux
    port map (
            O => \N__31504\,
            I => \N__31499\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__31499\,
            I => \N__31496\
        );

    \I__5711\ : Span4Mux_v
    port map (
            O => \N__31496\,
            I => \N__31492\
        );

    \I__5710\ : InMux
    port map (
            O => \N__31495\,
            I => \N__31489\
        );

    \I__5709\ : Span4Mux_v
    port map (
            O => \N__31492\,
            I => \N__31486\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__31489\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__5707\ : Odrv4
    port map (
            O => \N__31486\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__5706\ : InMux
    port map (
            O => \N__31481\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__5705\ : InMux
    port map (
            O => \N__31478\,
            I => \N__31475\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__31475\,
            I => \N__31471\
        );

    \I__5703\ : InMux
    port map (
            O => \N__31474\,
            I => \N__31468\
        );

    \I__5702\ : Span4Mux_h
    port map (
            O => \N__31471\,
            I => \N__31465\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__31468\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__5700\ : Odrv4
    port map (
            O => \N__31465\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__5699\ : InMux
    port map (
            O => \N__31460\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__5698\ : InMux
    port map (
            O => \N__31457\,
            I => \N__31454\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__31454\,
            I => \N__31450\
        );

    \I__5696\ : InMux
    port map (
            O => \N__31453\,
            I => \N__31447\
        );

    \I__5695\ : Span4Mux_v
    port map (
            O => \N__31450\,
            I => \N__31444\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__31447\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__31444\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__5692\ : InMux
    port map (
            O => \N__31439\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__5691\ : InMux
    port map (
            O => \N__31436\,
            I => \N__31433\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__31433\,
            I => \N__31429\
        );

    \I__5689\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31426\
        );

    \I__5688\ : Span4Mux_v
    port map (
            O => \N__31429\,
            I => \N__31423\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__31426\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__5686\ : Odrv4
    port map (
            O => \N__31423\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__5685\ : InMux
    port map (
            O => \N__31418\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__5684\ : InMux
    port map (
            O => \N__31415\,
            I => \N__31412\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__31412\,
            I => \N__31408\
        );

    \I__5682\ : InMux
    port map (
            O => \N__31411\,
            I => \N__31405\
        );

    \I__5681\ : Span4Mux_h
    port map (
            O => \N__31408\,
            I => \N__31402\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__31405\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__5679\ : Odrv4
    port map (
            O => \N__31402\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__5678\ : InMux
    port map (
            O => \N__31397\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__5677\ : InMux
    port map (
            O => \N__31394\,
            I => \N__31391\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__31391\,
            I => \N__31387\
        );

    \I__5675\ : InMux
    port map (
            O => \N__31390\,
            I => \N__31384\
        );

    \I__5674\ : Span4Mux_h
    port map (
            O => \N__31387\,
            I => \N__31381\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__31384\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__5672\ : Odrv4
    port map (
            O => \N__31381\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__5671\ : InMux
    port map (
            O => \N__31376\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__5670\ : InMux
    port map (
            O => \N__31373\,
            I => \N__31370\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__31370\,
            I => \N__31366\
        );

    \I__5668\ : InMux
    port map (
            O => \N__31369\,
            I => \N__31363\
        );

    \I__5667\ : Span4Mux_v
    port map (
            O => \N__31366\,
            I => \N__31360\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__31363\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__31360\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__5664\ : InMux
    port map (
            O => \N__31355\,
            I => \bfn_12_11_0_\
        );

    \I__5663\ : InMux
    port map (
            O => \N__31352\,
            I => \N__31349\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__31349\,
            I => \N__31345\
        );

    \I__5661\ : InMux
    port map (
            O => \N__31348\,
            I => \N__31342\
        );

    \I__5660\ : Span4Mux_v
    port map (
            O => \N__31345\,
            I => \N__31339\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__31342\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__5658\ : Odrv4
    port map (
            O => \N__31339\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__5657\ : InMux
    port map (
            O => \N__31334\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__5656\ : InMux
    port map (
            O => \N__31331\,
            I => \N__31328\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__31328\,
            I => \N__31324\
        );

    \I__5654\ : InMux
    port map (
            O => \N__31327\,
            I => \N__31321\
        );

    \I__5653\ : Span4Mux_h
    port map (
            O => \N__31324\,
            I => \N__31318\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__31321\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__5651\ : Odrv4
    port map (
            O => \N__31318\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__5650\ : InMux
    port map (
            O => \N__31313\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__5649\ : InMux
    port map (
            O => \N__31310\,
            I => \N__31306\
        );

    \I__5648\ : InMux
    port map (
            O => \N__31309\,
            I => \N__31302\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__31306\,
            I => \N__31299\
        );

    \I__5646\ : InMux
    port map (
            O => \N__31305\,
            I => \N__31296\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__31302\,
            I => \N__31289\
        );

    \I__5644\ : Span12Mux_v
    port map (
            O => \N__31299\,
            I => \N__31289\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__31296\,
            I => \N__31289\
        );

    \I__5642\ : Odrv12
    port map (
            O => \N__31289\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__5641\ : CascadeMux
    port map (
            O => \N__31286\,
            I => \N__31282\
        );

    \I__5640\ : CascadeMux
    port map (
            O => \N__31285\,
            I => \N__31279\
        );

    \I__5639\ : InMux
    port map (
            O => \N__31282\,
            I => \N__31276\
        );

    \I__5638\ : InMux
    port map (
            O => \N__31279\,
            I => \N__31273\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__31276\,
            I => \N__31270\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__31273\,
            I => \N__31267\
        );

    \I__5635\ : Span4Mux_v
    port map (
            O => \N__31270\,
            I => \N__31264\
        );

    \I__5634\ : Span4Mux_h
    port map (
            O => \N__31267\,
            I => \N__31261\
        );

    \I__5633\ : Odrv4
    port map (
            O => \N__31264\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\
        );

    \I__5632\ : Odrv4
    port map (
            O => \N__31261\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\
        );

    \I__5631\ : CascadeMux
    port map (
            O => \N__31256\,
            I => \N__31253\
        );

    \I__5630\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31250\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__31250\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\
        );

    \I__5628\ : InMux
    port map (
            O => \N__31247\,
            I => \N__31244\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__31244\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\
        );

    \I__5626\ : InMux
    port map (
            O => \N__31241\,
            I => \N__31238\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__31238\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\
        );

    \I__5624\ : InMux
    port map (
            O => \N__31235\,
            I => \N__31231\
        );

    \I__5623\ : CascadeMux
    port map (
            O => \N__31234\,
            I => \N__31228\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__31231\,
            I => \N__31225\
        );

    \I__5621\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31222\
        );

    \I__5620\ : Span4Mux_v
    port map (
            O => \N__31225\,
            I => \N__31219\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__31222\,
            I => \N__31214\
        );

    \I__5618\ : Span4Mux_h
    port map (
            O => \N__31219\,
            I => \N__31211\
        );

    \I__5617\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31208\
        );

    \I__5616\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31205\
        );

    \I__5615\ : Odrv12
    port map (
            O => \N__31214\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__5614\ : Odrv4
    port map (
            O => \N__31211\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__31208\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__31205\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__5611\ : InMux
    port map (
            O => \N__31196\,
            I => \N__31193\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__31193\,
            I => \N__31190\
        );

    \I__5609\ : Span4Mux_v
    port map (
            O => \N__31190\,
            I => \N__31186\
        );

    \I__5608\ : InMux
    port map (
            O => \N__31189\,
            I => \N__31183\
        );

    \I__5607\ : Odrv4
    port map (
            O => \N__31186\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__31183\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__5605\ : InMux
    port map (
            O => \N__31178\,
            I => \N__31175\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__31175\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\
        );

    \I__5603\ : InMux
    port map (
            O => \N__31172\,
            I => \N__31168\
        );

    \I__5602\ : InMux
    port map (
            O => \N__31171\,
            I => \N__31164\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__31168\,
            I => \N__31161\
        );

    \I__5600\ : CascadeMux
    port map (
            O => \N__31167\,
            I => \N__31158\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__31164\,
            I => \N__31155\
        );

    \I__5598\ : Span4Mux_v
    port map (
            O => \N__31161\,
            I => \N__31152\
        );

    \I__5597\ : InMux
    port map (
            O => \N__31158\,
            I => \N__31149\
        );

    \I__5596\ : Span12Mux_h
    port map (
            O => \N__31155\,
            I => \N__31146\
        );

    \I__5595\ : Span4Mux_h
    port map (
            O => \N__31152\,
            I => \N__31143\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__31149\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__5593\ : Odrv12
    port map (
            O => \N__31146\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__5592\ : Odrv4
    port map (
            O => \N__31143\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__5591\ : CascadeMux
    port map (
            O => \N__31136\,
            I => \N__31133\
        );

    \I__5590\ : InMux
    port map (
            O => \N__31133\,
            I => \N__31130\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__31130\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\
        );

    \I__5588\ : InMux
    port map (
            O => \N__31127\,
            I => \N__31124\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__31124\,
            I => \N__31120\
        );

    \I__5586\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31117\
        );

    \I__5585\ : Span4Mux_v
    port map (
            O => \N__31120\,
            I => \N__31114\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__31117\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__5583\ : Odrv4
    port map (
            O => \N__31114\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__5582\ : InMux
    port map (
            O => \N__31109\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__5581\ : InMux
    port map (
            O => \N__31106\,
            I => \N__31103\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__31103\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30\
        );

    \I__5579\ : InMux
    port map (
            O => \N__31100\,
            I => \N__31096\
        );

    \I__5578\ : CascadeMux
    port map (
            O => \N__31099\,
            I => \N__31093\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__31096\,
            I => \N__31090\
        );

    \I__5576\ : InMux
    port map (
            O => \N__31093\,
            I => \N__31087\
        );

    \I__5575\ : Span4Mux_h
    port map (
            O => \N__31090\,
            I => \N__31084\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__31087\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__31084\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__5572\ : InMux
    port map (
            O => \N__31079\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__5571\ : InMux
    port map (
            O => \N__31076\,
            I => \N__31073\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__31073\,
            I => \N__31068\
        );

    \I__5569\ : InMux
    port map (
            O => \N__31072\,
            I => \N__31065\
        );

    \I__5568\ : InMux
    port map (
            O => \N__31071\,
            I => \N__31062\
        );

    \I__5567\ : Span4Mux_v
    port map (
            O => \N__31068\,
            I => \N__31059\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__31065\,
            I => \N__31056\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__31062\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__5564\ : Odrv4
    port map (
            O => \N__31059\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__5563\ : Odrv4
    port map (
            O => \N__31056\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__5562\ : CascadeMux
    port map (
            O => \N__31049\,
            I => \N__31043\
        );

    \I__5561\ : InMux
    port map (
            O => \N__31048\,
            I => \N__31036\
        );

    \I__5560\ : InMux
    port map (
            O => \N__31047\,
            I => \N__31036\
        );

    \I__5559\ : InMux
    port map (
            O => \N__31046\,
            I => \N__31036\
        );

    \I__5558\ : InMux
    port map (
            O => \N__31043\,
            I => \N__31033\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__31036\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__31033\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5555\ : CascadeMux
    port map (
            O => \N__31028\,
            I => \N__31024\
        );

    \I__5554\ : InMux
    port map (
            O => \N__31027\,
            I => \N__31015\
        );

    \I__5553\ : InMux
    port map (
            O => \N__31024\,
            I => \N__31015\
        );

    \I__5552\ : InMux
    port map (
            O => \N__31023\,
            I => \N__31015\
        );

    \I__5551\ : InMux
    port map (
            O => \N__31022\,
            I => \N__31012\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__31015\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__31012\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__5548\ : IoInMux
    port map (
            O => \N__31007\,
            I => \N__31004\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__31004\,
            I => \N__31001\
        );

    \I__5546\ : IoSpan4Mux
    port map (
            O => \N__31001\,
            I => \N__30998\
        );

    \I__5545\ : Span4Mux_s0_v
    port map (
            O => \N__30998\,
            I => \N__30995\
        );

    \I__5544\ : Sp12to4
    port map (
            O => \N__30995\,
            I => \N__30992\
        );

    \I__5543\ : Span12Mux_v
    port map (
            O => \N__30992\,
            I => \N__30989\
        );

    \I__5542\ : Span12Mux_v
    port map (
            O => \N__30989\,
            I => \N__30985\
        );

    \I__5541\ : InMux
    port map (
            O => \N__30988\,
            I => \N__30982\
        );

    \I__5540\ : Odrv12
    port map (
            O => \N__30985\,
            I => test22_c
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__30982\,
            I => test22_c
        );

    \I__5538\ : InMux
    port map (
            O => \N__30977\,
            I => \N__30974\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__30974\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\
        );

    \I__5536\ : InMux
    port map (
            O => \N__30971\,
            I => \N__30968\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__30968\,
            I => \N__30964\
        );

    \I__5534\ : InMux
    port map (
            O => \N__30967\,
            I => \N__30961\
        );

    \I__5533\ : Span4Mux_s3_h
    port map (
            O => \N__30964\,
            I => \N__30958\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__30961\,
            I => \N__30955\
        );

    \I__5531\ : Span4Mux_v
    port map (
            O => \N__30958\,
            I => \N__30952\
        );

    \I__5530\ : Span12Mux_s8_h
    port map (
            O => \N__30955\,
            I => \N__30947\
        );

    \I__5529\ : Sp12to4
    port map (
            O => \N__30952\,
            I => \N__30947\
        );

    \I__5528\ : Odrv12
    port map (
            O => \N__30947\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__5527\ : InMux
    port map (
            O => \N__30944\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_22\
        );

    \I__5526\ : InMux
    port map (
            O => \N__30941\,
            I => \N__30938\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__30938\,
            I => \N__30935\
        );

    \I__5524\ : Span4Mux_v
    port map (
            O => \N__30935\,
            I => \N__30932\
        );

    \I__5523\ : Span4Mux_h
    port map (
            O => \N__30932\,
            I => \N__30929\
        );

    \I__5522\ : Span4Mux_h
    port map (
            O => \N__30929\,
            I => \N__30925\
        );

    \I__5521\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30922\
        );

    \I__5520\ : Span4Mux_h
    port map (
            O => \N__30925\,
            I => \N__30919\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__30922\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__5518\ : Odrv4
    port map (
            O => \N__30919\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__5517\ : InMux
    port map (
            O => \N__30914\,
            I => \bfn_11_22_0_\
        );

    \I__5516\ : InMux
    port map (
            O => \N__30911\,
            I => \N__30908\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__30908\,
            I => \N__30905\
        );

    \I__5514\ : Span4Mux_v
    port map (
            O => \N__30905\,
            I => \N__30902\
        );

    \I__5513\ : Span4Mux_h
    port map (
            O => \N__30902\,
            I => \N__30898\
        );

    \I__5512\ : InMux
    port map (
            O => \N__30901\,
            I => \N__30895\
        );

    \I__5511\ : Span4Mux_h
    port map (
            O => \N__30898\,
            I => \N__30892\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__30895\,
            I => \N__30887\
        );

    \I__5509\ : Span4Mux_h
    port map (
            O => \N__30892\,
            I => \N__30887\
        );

    \I__5508\ : Odrv4
    port map (
            O => \N__30887\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__5507\ : InMux
    port map (
            O => \N__30884\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_24\
        );

    \I__5506\ : InMux
    port map (
            O => \N__30881\,
            I => \N__30878\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__30878\,
            I => \N__30875\
        );

    \I__5504\ : Span4Mux_s1_h
    port map (
            O => \N__30875\,
            I => \N__30872\
        );

    \I__5503\ : Span4Mux_h
    port map (
            O => \N__30872\,
            I => \N__30868\
        );

    \I__5502\ : InMux
    port map (
            O => \N__30871\,
            I => \N__30865\
        );

    \I__5501\ : Span4Mux_h
    port map (
            O => \N__30868\,
            I => \N__30862\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__30865\,
            I => \N__30859\
        );

    \I__5499\ : Span4Mux_h
    port map (
            O => \N__30862\,
            I => \N__30856\
        );

    \I__5498\ : Odrv4
    port map (
            O => \N__30859\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__30856\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__5496\ : InMux
    port map (
            O => \N__30851\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_25\
        );

    \I__5495\ : InMux
    port map (
            O => \N__30848\,
            I => \N__30845\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__30845\,
            I => \N__30841\
        );

    \I__5493\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30838\
        );

    \I__5492\ : Span12Mux_s2_h
    port map (
            O => \N__30841\,
            I => \N__30835\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__30838\,
            I => \N__30832\
        );

    \I__5490\ : Span12Mux_h
    port map (
            O => \N__30835\,
            I => \N__30829\
        );

    \I__5489\ : Odrv4
    port map (
            O => \N__30832\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_27\
        );

    \I__5488\ : Odrv12
    port map (
            O => \N__30829\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_27\
        );

    \I__5487\ : InMux
    port map (
            O => \N__30824\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_26\
        );

    \I__5486\ : InMux
    port map (
            O => \N__30821\,
            I => \N__30818\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__30818\,
            I => \N__30815\
        );

    \I__5484\ : Span4Mux_s1_h
    port map (
            O => \N__30815\,
            I => \N__30812\
        );

    \I__5483\ : Span4Mux_h
    port map (
            O => \N__30812\,
            I => \N__30809\
        );

    \I__5482\ : Span4Mux_h
    port map (
            O => \N__30809\,
            I => \N__30805\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30808\,
            I => \N__30802\
        );

    \I__5480\ : Span4Mux_h
    port map (
            O => \N__30805\,
            I => \N__30799\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__30802\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__5478\ : Odrv4
    port map (
            O => \N__30799\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__5477\ : InMux
    port map (
            O => \N__30794\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_27\
        );

    \I__5476\ : InMux
    port map (
            O => \N__30791\,
            I => \N__30788\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__30788\,
            I => \N__30785\
        );

    \I__5474\ : Span4Mux_s3_h
    port map (
            O => \N__30785\,
            I => \N__30781\
        );

    \I__5473\ : InMux
    port map (
            O => \N__30784\,
            I => \N__30778\
        );

    \I__5472\ : Sp12to4
    port map (
            O => \N__30781\,
            I => \N__30775\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__30778\,
            I => \N__30770\
        );

    \I__5470\ : Span12Mux_s8_v
    port map (
            O => \N__30775\,
            I => \N__30770\
        );

    \I__5469\ : Odrv12
    port map (
            O => \N__30770\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__5468\ : InMux
    port map (
            O => \N__30767\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_28\
        );

    \I__5467\ : InMux
    port map (
            O => \N__30764\,
            I => \N__30761\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__30761\,
            I => \N__30758\
        );

    \I__5465\ : Span12Mux_s8_v
    port map (
            O => \N__30758\,
            I => \N__30754\
        );

    \I__5464\ : InMux
    port map (
            O => \N__30757\,
            I => \N__30751\
        );

    \I__5463\ : Span12Mux_h
    port map (
            O => \N__30754\,
            I => \N__30748\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__30751\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__5461\ : Odrv12
    port map (
            O => \N__30748\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__5460\ : InMux
    port map (
            O => \N__30743\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_29\
        );

    \I__5459\ : InMux
    port map (
            O => \N__30740\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_30\
        );

    \I__5458\ : InMux
    port map (
            O => \N__30737\,
            I => \N__30734\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__30734\,
            I => \N__30731\
        );

    \I__5456\ : Odrv4
    port map (
            O => \N__30731\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_31\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30725\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__30725\,
            I => \N__30722\
        );

    \I__5453\ : Span4Mux_v
    port map (
            O => \N__30722\,
            I => \N__30718\
        );

    \I__5452\ : InMux
    port map (
            O => \N__30721\,
            I => \N__30715\
        );

    \I__5451\ : Sp12to4
    port map (
            O => \N__30718\,
            I => \N__30712\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__30715\,
            I => \N__30709\
        );

    \I__5449\ : Span12Mux_h
    port map (
            O => \N__30712\,
            I => \N__30706\
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__30709\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__5447\ : Odrv12
    port map (
            O => \N__30706\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__5446\ : InMux
    port map (
            O => \N__30701\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_14\
        );

    \I__5445\ : InMux
    port map (
            O => \N__30698\,
            I => \N__30695\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__30695\,
            I => \N__30692\
        );

    \I__5443\ : Span4Mux_s2_h
    port map (
            O => \N__30692\,
            I => \N__30688\
        );

    \I__5442\ : InMux
    port map (
            O => \N__30691\,
            I => \N__30685\
        );

    \I__5441\ : Span4Mux_h
    port map (
            O => \N__30688\,
            I => \N__30682\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__30685\,
            I => \N__30679\
        );

    \I__5439\ : Span4Mux_h
    port map (
            O => \N__30682\,
            I => \N__30676\
        );

    \I__5438\ : Span4Mux_v
    port map (
            O => \N__30679\,
            I => \N__30673\
        );

    \I__5437\ : Span4Mux_v
    port map (
            O => \N__30676\,
            I => \N__30670\
        );

    \I__5436\ : Odrv4
    port map (
            O => \N__30673\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__5435\ : Odrv4
    port map (
            O => \N__30670\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__5434\ : InMux
    port map (
            O => \N__30665\,
            I => \bfn_11_21_0_\
        );

    \I__5433\ : InMux
    port map (
            O => \N__30662\,
            I => \N__30659\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__30659\,
            I => \N__30656\
        );

    \I__5431\ : Span4Mux_v
    port map (
            O => \N__30656\,
            I => \N__30652\
        );

    \I__5430\ : InMux
    port map (
            O => \N__30655\,
            I => \N__30649\
        );

    \I__5429\ : Sp12to4
    port map (
            O => \N__30652\,
            I => \N__30646\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__30649\,
            I => \N__30643\
        );

    \I__5427\ : Span12Mux_h
    port map (
            O => \N__30646\,
            I => \N__30640\
        );

    \I__5426\ : Odrv12
    port map (
            O => \N__30643\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__5425\ : Odrv12
    port map (
            O => \N__30640\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__5424\ : InMux
    port map (
            O => \N__30635\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_16\
        );

    \I__5423\ : InMux
    port map (
            O => \N__30632\,
            I => \N__30629\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__30629\,
            I => \N__30626\
        );

    \I__5421\ : Span4Mux_s2_h
    port map (
            O => \N__30626\,
            I => \N__30623\
        );

    \I__5420\ : Span4Mux_h
    port map (
            O => \N__30623\,
            I => \N__30619\
        );

    \I__5419\ : InMux
    port map (
            O => \N__30622\,
            I => \N__30616\
        );

    \I__5418\ : Span4Mux_h
    port map (
            O => \N__30619\,
            I => \N__30613\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__30616\,
            I => \N__30610\
        );

    \I__5416\ : Span4Mux_v
    port map (
            O => \N__30613\,
            I => \N__30607\
        );

    \I__5415\ : Odrv4
    port map (
            O => \N__30610\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__5414\ : Odrv4
    port map (
            O => \N__30607\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__5413\ : InMux
    port map (
            O => \N__30602\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_17\
        );

    \I__5412\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30596\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__30596\,
            I => \N__30593\
        );

    \I__5410\ : Span4Mux_v
    port map (
            O => \N__30593\,
            I => \N__30589\
        );

    \I__5409\ : InMux
    port map (
            O => \N__30592\,
            I => \N__30586\
        );

    \I__5408\ : Sp12to4
    port map (
            O => \N__30589\,
            I => \N__30583\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__30586\,
            I => \N__30580\
        );

    \I__5406\ : Span12Mux_h
    port map (
            O => \N__30583\,
            I => \N__30577\
        );

    \I__5405\ : Odrv12
    port map (
            O => \N__30580\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__5404\ : Odrv12
    port map (
            O => \N__30577\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__5403\ : InMux
    port map (
            O => \N__30572\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_18\
        );

    \I__5402\ : InMux
    port map (
            O => \N__30569\,
            I => \N__30566\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__30566\,
            I => \N__30562\
        );

    \I__5400\ : InMux
    port map (
            O => \N__30565\,
            I => \N__30559\
        );

    \I__5399\ : Span12Mux_s2_h
    port map (
            O => \N__30562\,
            I => \N__30556\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__30559\,
            I => \N__30553\
        );

    \I__5397\ : Span12Mux_h
    port map (
            O => \N__30556\,
            I => \N__30550\
        );

    \I__5396\ : Odrv4
    port map (
            O => \N__30553\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__5395\ : Odrv12
    port map (
            O => \N__30550\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__5394\ : InMux
    port map (
            O => \N__30545\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_19\
        );

    \I__5393\ : InMux
    port map (
            O => \N__30542\,
            I => \N__30539\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__30539\,
            I => \N__30536\
        );

    \I__5391\ : Span4Mux_s1_h
    port map (
            O => \N__30536\,
            I => \N__30532\
        );

    \I__5390\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30529\
        );

    \I__5389\ : Span4Mux_v
    port map (
            O => \N__30532\,
            I => \N__30526\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__30529\,
            I => \N__30523\
        );

    \I__5387\ : Sp12to4
    port map (
            O => \N__30526\,
            I => \N__30520\
        );

    \I__5386\ : Odrv4
    port map (
            O => \N__30523\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__5385\ : Odrv12
    port map (
            O => \N__30520\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__5384\ : InMux
    port map (
            O => \N__30515\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_20\
        );

    \I__5383\ : InMux
    port map (
            O => \N__30512\,
            I => \N__30509\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__30509\,
            I => \N__30505\
        );

    \I__5381\ : InMux
    port map (
            O => \N__30508\,
            I => \N__30502\
        );

    \I__5380\ : Span12Mux_s9_v
    port map (
            O => \N__30505\,
            I => \N__30499\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__30502\,
            I => \N__30494\
        );

    \I__5378\ : Span12Mux_h
    port map (
            O => \N__30499\,
            I => \N__30494\
        );

    \I__5377\ : Odrv12
    port map (
            O => \N__30494\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__5376\ : InMux
    port map (
            O => \N__30491\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_21\
        );

    \I__5375\ : InMux
    port map (
            O => \N__30488\,
            I => \N__30485\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__30485\,
            I => \N__30482\
        );

    \I__5373\ : Span4Mux_s3_h
    port map (
            O => \N__30482\,
            I => \N__30478\
        );

    \I__5372\ : InMux
    port map (
            O => \N__30481\,
            I => \N__30475\
        );

    \I__5371\ : Span4Mux_h
    port map (
            O => \N__30478\,
            I => \N__30472\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__30475\,
            I => \N__30469\
        );

    \I__5369\ : Span4Mux_h
    port map (
            O => \N__30472\,
            I => \N__30466\
        );

    \I__5368\ : Span12Mux_s9_h
    port map (
            O => \N__30469\,
            I => \N__30463\
        );

    \I__5367\ : Span4Mux_v
    port map (
            O => \N__30466\,
            I => \N__30460\
        );

    \I__5366\ : Odrv12
    port map (
            O => \N__30463\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__5365\ : Odrv4
    port map (
            O => \N__30460\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__5364\ : InMux
    port map (
            O => \N__30455\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__5363\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30449\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__30449\,
            I => \N__30445\
        );

    \I__5361\ : InMux
    port map (
            O => \N__30448\,
            I => \N__30442\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__30445\,
            I => \N__30439\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__30442\,
            I => \N__30436\
        );

    \I__5358\ : Span4Mux_h
    port map (
            O => \N__30439\,
            I => \N__30433\
        );

    \I__5357\ : Span12Mux_v
    port map (
            O => \N__30436\,
            I => \N__30430\
        );

    \I__5356\ : Odrv4
    port map (
            O => \N__30433\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__5355\ : Odrv12
    port map (
            O => \N__30430\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__5354\ : InMux
    port map (
            O => \N__30425\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__5353\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30418\
        );

    \I__5352\ : InMux
    port map (
            O => \N__30421\,
            I => \N__30415\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__30418\,
            I => \N__30412\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__30415\,
            I => \N__30409\
        );

    \I__5349\ : Span4Mux_h
    port map (
            O => \N__30412\,
            I => \N__30406\
        );

    \I__5348\ : Span4Mux_v
    port map (
            O => \N__30409\,
            I => \N__30401\
        );

    \I__5347\ : Span4Mux_v
    port map (
            O => \N__30406\,
            I => \N__30401\
        );

    \I__5346\ : Sp12to4
    port map (
            O => \N__30401\,
            I => \N__30398\
        );

    \I__5345\ : Span12Mux_s11_h
    port map (
            O => \N__30398\,
            I => \N__30395\
        );

    \I__5344\ : Odrv12
    port map (
            O => \N__30395\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__5343\ : InMux
    port map (
            O => \N__30392\,
            I => \bfn_11_20_0_\
        );

    \I__5342\ : InMux
    port map (
            O => \N__30389\,
            I => \N__30386\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__30386\,
            I => \N__30383\
        );

    \I__5340\ : Span4Mux_v
    port map (
            O => \N__30383\,
            I => \N__30380\
        );

    \I__5339\ : Sp12to4
    port map (
            O => \N__30380\,
            I => \N__30376\
        );

    \I__5338\ : InMux
    port map (
            O => \N__30379\,
            I => \N__30373\
        );

    \I__5337\ : Span12Mux_s6_h
    port map (
            O => \N__30376\,
            I => \N__30370\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__30373\,
            I => \N__30365\
        );

    \I__5335\ : Span12Mux_v
    port map (
            O => \N__30370\,
            I => \N__30365\
        );

    \I__5334\ : Odrv12
    port map (
            O => \N__30365\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__5333\ : InMux
    port map (
            O => \N__30362\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__5332\ : InMux
    port map (
            O => \N__30359\,
            I => \N__30356\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__30356\,
            I => \N__30353\
        );

    \I__5330\ : Span4Mux_v
    port map (
            O => \N__30353\,
            I => \N__30349\
        );

    \I__5329\ : InMux
    port map (
            O => \N__30352\,
            I => \N__30346\
        );

    \I__5328\ : Sp12to4
    port map (
            O => \N__30349\,
            I => \N__30343\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__30346\,
            I => \N__30340\
        );

    \I__5326\ : Span12Mux_s11_h
    port map (
            O => \N__30343\,
            I => \N__30337\
        );

    \I__5325\ : Odrv12
    port map (
            O => \N__30340\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__5324\ : Odrv12
    port map (
            O => \N__30337\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__5323\ : InMux
    port map (
            O => \N__30332\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__5322\ : InMux
    port map (
            O => \N__30329\,
            I => \N__30326\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__30326\,
            I => \N__30323\
        );

    \I__5320\ : Span4Mux_v
    port map (
            O => \N__30323\,
            I => \N__30319\
        );

    \I__5319\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30316\
        );

    \I__5318\ : Sp12to4
    port map (
            O => \N__30319\,
            I => \N__30313\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__30316\,
            I => \N__30310\
        );

    \I__5316\ : Span12Mux_s11_h
    port map (
            O => \N__30313\,
            I => \N__30307\
        );

    \I__5315\ : Odrv12
    port map (
            O => \N__30310\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__5314\ : Odrv12
    port map (
            O => \N__30307\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__5313\ : InMux
    port map (
            O => \N__30302\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__5312\ : InMux
    port map (
            O => \N__30299\,
            I => \N__30295\
        );

    \I__5311\ : InMux
    port map (
            O => \N__30298\,
            I => \N__30292\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__30295\,
            I => \N__30289\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__30292\,
            I => \N__30286\
        );

    \I__5308\ : Span12Mux_s11_h
    port map (
            O => \N__30289\,
            I => \N__30283\
        );

    \I__5307\ : Odrv12
    port map (
            O => \N__30286\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__5306\ : Odrv12
    port map (
            O => \N__30283\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__5305\ : InMux
    port map (
            O => \N__30278\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__5304\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30272\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__30272\,
            I => \N__30269\
        );

    \I__5302\ : Span4Mux_s3_h
    port map (
            O => \N__30269\,
            I => \N__30265\
        );

    \I__5301\ : InMux
    port map (
            O => \N__30268\,
            I => \N__30262\
        );

    \I__5300\ : Span4Mux_v
    port map (
            O => \N__30265\,
            I => \N__30259\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__30262\,
            I => \N__30256\
        );

    \I__5298\ : Span4Mux_h
    port map (
            O => \N__30259\,
            I => \N__30253\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__30256\,
            I => \N__30248\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__30253\,
            I => \N__30248\
        );

    \I__5295\ : Odrv4
    port map (
            O => \N__30248\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__5294\ : InMux
    port map (
            O => \N__30245\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__5293\ : InMux
    port map (
            O => \N__30242\,
            I => \N__30239\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__30239\,
            I => \N__30236\
        );

    \I__5291\ : Span4Mux_v
    port map (
            O => \N__30236\,
            I => \N__30232\
        );

    \I__5290\ : InMux
    port map (
            O => \N__30235\,
            I => \N__30229\
        );

    \I__5289\ : Sp12to4
    port map (
            O => \N__30232\,
            I => \N__30226\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__30229\,
            I => \N__30223\
        );

    \I__5287\ : Span12Mux_s11_h
    port map (
            O => \N__30226\,
            I => \N__30220\
        );

    \I__5286\ : Odrv12
    port map (
            O => \N__30223\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__5285\ : Odrv12
    port map (
            O => \N__30220\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__5284\ : InMux
    port map (
            O => \N__30215\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__5283\ : InMux
    port map (
            O => \N__30212\,
            I => \N__30209\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__30209\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__5281\ : InMux
    port map (
            O => \N__30206\,
            I => \N__30203\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__30203\,
            I => \N__30200\
        );

    \I__5279\ : Span4Mux_s3_h
    port map (
            O => \N__30200\,
            I => \N__30196\
        );

    \I__5278\ : InMux
    port map (
            O => \N__30199\,
            I => \N__30193\
        );

    \I__5277\ : Span4Mux_v
    port map (
            O => \N__30196\,
            I => \N__30190\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__30193\,
            I => \N__30187\
        );

    \I__5275\ : Span4Mux_h
    port map (
            O => \N__30190\,
            I => \N__30184\
        );

    \I__5274\ : Span12Mux_s6_h
    port map (
            O => \N__30187\,
            I => \N__30181\
        );

    \I__5273\ : Span4Mux_h
    port map (
            O => \N__30184\,
            I => \N__30178\
        );

    \I__5272\ : Odrv12
    port map (
            O => \N__30181\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__5271\ : Odrv4
    port map (
            O => \N__30178\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__5270\ : InMux
    port map (
            O => \N__30173\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__5269\ : InMux
    port map (
            O => \N__30170\,
            I => \N__30167\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__30167\,
            I => \N__30163\
        );

    \I__5267\ : InMux
    port map (
            O => \N__30166\,
            I => \N__30160\
        );

    \I__5266\ : Span4Mux_v
    port map (
            O => \N__30163\,
            I => \N__30157\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__30160\,
            I => \N__30154\
        );

    \I__5264\ : Sp12to4
    port map (
            O => \N__30157\,
            I => \N__30151\
        );

    \I__5263\ : Span12Mux_v
    port map (
            O => \N__30154\,
            I => \N__30148\
        );

    \I__5262\ : Span12Mux_s11_h
    port map (
            O => \N__30151\,
            I => \N__30145\
        );

    \I__5261\ : Odrv12
    port map (
            O => \N__30148\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__5260\ : Odrv12
    port map (
            O => \N__30145\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__5259\ : InMux
    port map (
            O => \N__30140\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__5258\ : InMux
    port map (
            O => \N__30137\,
            I => \N__30134\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__30134\,
            I => \N__30130\
        );

    \I__5256\ : InMux
    port map (
            O => \N__30133\,
            I => \N__30127\
        );

    \I__5255\ : Span4Mux_h
    port map (
            O => \N__30130\,
            I => \N__30124\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__30127\,
            I => \N__30121\
        );

    \I__5253\ : Sp12to4
    port map (
            O => \N__30124\,
            I => \N__30118\
        );

    \I__5252\ : Span12Mux_s4_h
    port map (
            O => \N__30121\,
            I => \N__30113\
        );

    \I__5251\ : Span12Mux_v
    port map (
            O => \N__30118\,
            I => \N__30113\
        );

    \I__5250\ : Odrv12
    port map (
            O => \N__30113\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__5249\ : InMux
    port map (
            O => \N__30110\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__5248\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30103\
        );

    \I__5247\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30100\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__30103\,
            I => \N__30097\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__30100\,
            I => \N__30094\
        );

    \I__5244\ : Span4Mux_v
    port map (
            O => \N__30097\,
            I => \N__30091\
        );

    \I__5243\ : Span4Mux_h
    port map (
            O => \N__30094\,
            I => \N__30088\
        );

    \I__5242\ : Sp12to4
    port map (
            O => \N__30091\,
            I => \N__30085\
        );

    \I__5241\ : Span4Mux_h
    port map (
            O => \N__30088\,
            I => \N__30082\
        );

    \I__5240\ : Span12Mux_s11_h
    port map (
            O => \N__30085\,
            I => \N__30079\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__30082\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__5238\ : Odrv12
    port map (
            O => \N__30079\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__5237\ : InMux
    port map (
            O => \N__30074\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__5236\ : InMux
    port map (
            O => \N__30071\,
            I => \N__30067\
        );

    \I__5235\ : InMux
    port map (
            O => \N__30070\,
            I => \N__30064\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__30067\,
            I => \N__30061\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__30064\,
            I => \N__30058\
        );

    \I__5232\ : Span4Mux_s2_h
    port map (
            O => \N__30061\,
            I => \N__30055\
        );

    \I__5231\ : Span4Mux_v
    port map (
            O => \N__30058\,
            I => \N__30052\
        );

    \I__5230\ : Sp12to4
    port map (
            O => \N__30055\,
            I => \N__30049\
        );

    \I__5229\ : Sp12to4
    port map (
            O => \N__30052\,
            I => \N__30044\
        );

    \I__5228\ : Span12Mux_v
    port map (
            O => \N__30049\,
            I => \N__30044\
        );

    \I__5227\ : Odrv12
    port map (
            O => \N__30044\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__5226\ : InMux
    port map (
            O => \N__30041\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__30038\,
            I => \N__30034\
        );

    \I__5224\ : InMux
    port map (
            O => \N__30037\,
            I => \N__30028\
        );

    \I__5223\ : InMux
    port map (
            O => \N__30034\,
            I => \N__30028\
        );

    \I__5222\ : InMux
    port map (
            O => \N__30033\,
            I => \N__30025\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__30028\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__30025\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__5219\ : InMux
    port map (
            O => \N__30020\,
            I => \N__30016\
        );

    \I__5218\ : InMux
    port map (
            O => \N__30019\,
            I => \N__30013\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__30016\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__30013\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__5215\ : InMux
    port map (
            O => \N__30008\,
            I => \N__30004\
        );

    \I__5214\ : InMux
    port map (
            O => \N__30007\,
            I => \N__30001\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__30004\,
            I => \N__29996\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__30001\,
            I => \N__29996\
        );

    \I__5211\ : Span4Mux_s3_v
    port map (
            O => \N__29996\,
            I => \N__29991\
        );

    \I__5210\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29988\
        );

    \I__5209\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29985\
        );

    \I__5208\ : Span4Mux_h
    port map (
            O => \N__29991\,
            I => \N__29982\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__29988\,
            I => \N__29979\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__29985\,
            I => \N__29976\
        );

    \I__5205\ : Sp12to4
    port map (
            O => \N__29982\,
            I => \N__29973\
        );

    \I__5204\ : Span4Mux_h
    port map (
            O => \N__29979\,
            I => \N__29970\
        );

    \I__5203\ : Span4Mux_v
    port map (
            O => \N__29976\,
            I => \N__29967\
        );

    \I__5202\ : Span12Mux_s11_v
    port map (
            O => \N__29973\,
            I => \N__29962\
        );

    \I__5201\ : Sp12to4
    port map (
            O => \N__29970\,
            I => \N__29962\
        );

    \I__5200\ : Span4Mux_v
    port map (
            O => \N__29967\,
            I => \N__29959\
        );

    \I__5199\ : Span12Mux_v
    port map (
            O => \N__29962\,
            I => \N__29956\
        );

    \I__5198\ : Sp12to4
    port map (
            O => \N__29959\,
            I => \N__29953\
        );

    \I__5197\ : Span12Mux_h
    port map (
            O => \N__29956\,
            I => \N__29950\
        );

    \I__5196\ : Span12Mux_h
    port map (
            O => \N__29953\,
            I => \N__29947\
        );

    \I__5195\ : Odrv12
    port map (
            O => \N__29950\,
            I => start_stop_c
        );

    \I__5194\ : Odrv12
    port map (
            O => \N__29947\,
            I => start_stop_c
        );

    \I__5193\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29939\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__29939\,
            I => \N__29936\
        );

    \I__5191\ : Span4Mux_v
    port map (
            O => \N__29936\,
            I => \N__29931\
        );

    \I__5190\ : InMux
    port map (
            O => \N__29935\,
            I => \N__29928\
        );

    \I__5189\ : InMux
    port map (
            O => \N__29934\,
            I => \N__29925\
        );

    \I__5188\ : Sp12to4
    port map (
            O => \N__29931\,
            I => \N__29918\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__29928\,
            I => \N__29918\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__29925\,
            I => \N__29918\
        );

    \I__5185\ : Span12Mux_h
    port map (
            O => \N__29918\,
            I => \N__29915\
        );

    \I__5184\ : Span12Mux_v
    port map (
            O => \N__29915\,
            I => \N__29912\
        );

    \I__5183\ : Odrv12
    port map (
            O => \N__29912\,
            I => il_max_comp2_c
        );

    \I__5182\ : CascadeMux
    port map (
            O => \N__29909\,
            I => \phase_controller_inst1_N_54_cascade_\
        );

    \I__5181\ : InMux
    port map (
            O => \N__29906\,
            I => \N__29903\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__29903\,
            I => \N__29899\
        );

    \I__5179\ : InMux
    port map (
            O => \N__29902\,
            I => \N__29896\
        );

    \I__5178\ : Odrv4
    port map (
            O => \N__29899\,
            I => \phase_controller_inst2.N_54\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__29896\,
            I => \phase_controller_inst2.N_54\
        );

    \I__5176\ : CascadeMux
    port map (
            O => \N__29891\,
            I => \N__29888\
        );

    \I__5175\ : InMux
    port map (
            O => \N__29888\,
            I => \N__29884\
        );

    \I__5174\ : InMux
    port map (
            O => \N__29887\,
            I => \N__29881\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__29884\,
            I => \N__29875\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__29881\,
            I => \N__29875\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29880\,
            I => \N__29871\
        );

    \I__5170\ : Span12Mux_v
    port map (
            O => \N__29875\,
            I => \N__29868\
        );

    \I__5169\ : InMux
    port map (
            O => \N__29874\,
            I => \N__29865\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__29871\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__5167\ : Odrv12
    port map (
            O => \N__29868\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__29865\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__5165\ : CEMux
    port map (
            O => \N__29858\,
            I => \N__29853\
        );

    \I__5164\ : CEMux
    port map (
            O => \N__29857\,
            I => \N__29849\
        );

    \I__5163\ : CEMux
    port map (
            O => \N__29856\,
            I => \N__29846\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__29853\,
            I => \N__29843\
        );

    \I__5161\ : CEMux
    port map (
            O => \N__29852\,
            I => \N__29840\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__29849\,
            I => \N__29837\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__29846\,
            I => \N__29834\
        );

    \I__5158\ : Span4Mux_v
    port map (
            O => \N__29843\,
            I => \N__29829\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__29840\,
            I => \N__29829\
        );

    \I__5156\ : Span4Mux_v
    port map (
            O => \N__29837\,
            I => \N__29826\
        );

    \I__5155\ : Span4Mux_v
    port map (
            O => \N__29834\,
            I => \N__29823\
        );

    \I__5154\ : Span4Mux_h
    port map (
            O => \N__29829\,
            I => \N__29820\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__29826\,
            I => \delay_measurement_inst.delay_tr_timer.N_166_i\
        );

    \I__5152\ : Odrv4
    port map (
            O => \N__29823\,
            I => \delay_measurement_inst.delay_tr_timer.N_166_i\
        );

    \I__5151\ : Odrv4
    port map (
            O => \N__29820\,
            I => \delay_measurement_inst.delay_tr_timer.N_166_i\
        );

    \I__5150\ : CascadeMux
    port map (
            O => \N__29813\,
            I => \N__29809\
        );

    \I__5149\ : InMux
    port map (
            O => \N__29812\,
            I => \N__29804\
        );

    \I__5148\ : InMux
    port map (
            O => \N__29809\,
            I => \N__29799\
        );

    \I__5147\ : InMux
    port map (
            O => \N__29808\,
            I => \N__29799\
        );

    \I__5146\ : InMux
    port map (
            O => \N__29807\,
            I => \N__29796\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__29804\,
            I => \N__29793\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__29799\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__29796\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__29793\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5141\ : InMux
    port map (
            O => \N__29786\,
            I => \N__29780\
        );

    \I__5140\ : InMux
    port map (
            O => \N__29785\,
            I => \N__29777\
        );

    \I__5139\ : InMux
    port map (
            O => \N__29784\,
            I => \N__29772\
        );

    \I__5138\ : InMux
    port map (
            O => \N__29783\,
            I => \N__29772\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__29780\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__29777\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__29772\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__5134\ : InMux
    port map (
            O => \N__29765\,
            I => \N__29753\
        );

    \I__5133\ : InMux
    port map (
            O => \N__29764\,
            I => \N__29753\
        );

    \I__5132\ : InMux
    port map (
            O => \N__29763\,
            I => \N__29753\
        );

    \I__5131\ : InMux
    port map (
            O => \N__29762\,
            I => \N__29753\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__29753\,
            I => \N__29728\
        );

    \I__5129\ : InMux
    port map (
            O => \N__29752\,
            I => \N__29719\
        );

    \I__5128\ : InMux
    port map (
            O => \N__29751\,
            I => \N__29719\
        );

    \I__5127\ : InMux
    port map (
            O => \N__29750\,
            I => \N__29719\
        );

    \I__5126\ : InMux
    port map (
            O => \N__29749\,
            I => \N__29719\
        );

    \I__5125\ : InMux
    port map (
            O => \N__29748\,
            I => \N__29710\
        );

    \I__5124\ : InMux
    port map (
            O => \N__29747\,
            I => \N__29710\
        );

    \I__5123\ : InMux
    port map (
            O => \N__29746\,
            I => \N__29710\
        );

    \I__5122\ : InMux
    port map (
            O => \N__29745\,
            I => \N__29710\
        );

    \I__5121\ : InMux
    port map (
            O => \N__29744\,
            I => \N__29701\
        );

    \I__5120\ : InMux
    port map (
            O => \N__29743\,
            I => \N__29701\
        );

    \I__5119\ : InMux
    port map (
            O => \N__29742\,
            I => \N__29692\
        );

    \I__5118\ : InMux
    port map (
            O => \N__29741\,
            I => \N__29692\
        );

    \I__5117\ : InMux
    port map (
            O => \N__29740\,
            I => \N__29692\
        );

    \I__5116\ : InMux
    port map (
            O => \N__29739\,
            I => \N__29692\
        );

    \I__5115\ : InMux
    port map (
            O => \N__29738\,
            I => \N__29683\
        );

    \I__5114\ : InMux
    port map (
            O => \N__29737\,
            I => \N__29683\
        );

    \I__5113\ : InMux
    port map (
            O => \N__29736\,
            I => \N__29683\
        );

    \I__5112\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29683\
        );

    \I__5111\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29674\
        );

    \I__5110\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29674\
        );

    \I__5109\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29674\
        );

    \I__5108\ : InMux
    port map (
            O => \N__29731\,
            I => \N__29674\
        );

    \I__5107\ : Span4Mux_v
    port map (
            O => \N__29728\,
            I => \N__29667\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__29719\,
            I => \N__29667\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__29710\,
            I => \N__29667\
        );

    \I__5104\ : InMux
    port map (
            O => \N__29709\,
            I => \N__29658\
        );

    \I__5103\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29658\
        );

    \I__5102\ : InMux
    port map (
            O => \N__29707\,
            I => \N__29658\
        );

    \I__5101\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29658\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__29701\,
            I => \N__29645\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__29692\,
            I => \N__29645\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__29683\,
            I => \N__29645\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__29674\,
            I => \N__29645\
        );

    \I__5096\ : Span4Mux_h
    port map (
            O => \N__29667\,
            I => \N__29645\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__29658\,
            I => \N__29645\
        );

    \I__5094\ : Span4Mux_v
    port map (
            O => \N__29645\,
            I => \N__29642\
        );

    \I__5093\ : Odrv4
    port map (
            O => \N__29642\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__5092\ : CascadeMux
    port map (
            O => \N__29639\,
            I => \current_shift_inst.control_input_axb_0_cascade_\
        );

    \I__5091\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29633\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__29633\,
            I => \N__29629\
        );

    \I__5089\ : InMux
    port map (
            O => \N__29632\,
            I => \N__29626\
        );

    \I__5088\ : Span4Mux_v
    port map (
            O => \N__29629\,
            I => \N__29623\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__29626\,
            I => \N__29620\
        );

    \I__5086\ : Sp12to4
    port map (
            O => \N__29623\,
            I => \N__29617\
        );

    \I__5085\ : Span4Mux_h
    port map (
            O => \N__29620\,
            I => \N__29614\
        );

    \I__5084\ : Span12Mux_s11_h
    port map (
            O => \N__29617\,
            I => \N__29611\
        );

    \I__5083\ : Odrv4
    port map (
            O => \N__29614\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__5082\ : Odrv12
    port map (
            O => \N__29611\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__5081\ : InMux
    port map (
            O => \N__29606\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__5080\ : InMux
    port map (
            O => \N__29603\,
            I => \bfn_11_14_0_\
        );

    \I__5079\ : InMux
    port map (
            O => \N__29600\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__5078\ : InMux
    port map (
            O => \N__29597\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__5077\ : InMux
    port map (
            O => \N__29594\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__5076\ : InMux
    port map (
            O => \N__29591\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__5075\ : InMux
    port map (
            O => \N__29588\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__5074\ : InMux
    port map (
            O => \N__29585\,
            I => \N__29581\
        );

    \I__5073\ : InMux
    port map (
            O => \N__29584\,
            I => \N__29578\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__29581\,
            I => \N__29572\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__29578\,
            I => \N__29572\
        );

    \I__5070\ : InMux
    port map (
            O => \N__29577\,
            I => \N__29567\
        );

    \I__5069\ : Span4Mux_v
    port map (
            O => \N__29572\,
            I => \N__29564\
        );

    \I__5068\ : InMux
    port map (
            O => \N__29571\,
            I => \N__29559\
        );

    \I__5067\ : InMux
    port map (
            O => \N__29570\,
            I => \N__29559\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__29567\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__5065\ : Odrv4
    port map (
            O => \N__29564\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__29559\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__5063\ : InMux
    port map (
            O => \N__29552\,
            I => \N__29549\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__29549\,
            I => \N__29545\
        );

    \I__5061\ : InMux
    port map (
            O => \N__29548\,
            I => \N__29541\
        );

    \I__5060\ : Span4Mux_v
    port map (
            O => \N__29545\,
            I => \N__29538\
        );

    \I__5059\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29535\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__29541\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__5057\ : Odrv4
    port map (
            O => \N__29538\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__29535\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__5055\ : InMux
    port map (
            O => \N__29528\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__5054\ : InMux
    port map (
            O => \N__29525\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__5053\ : InMux
    port map (
            O => \N__29522\,
            I => \bfn_11_13_0_\
        );

    \I__5052\ : InMux
    port map (
            O => \N__29519\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__5051\ : InMux
    port map (
            O => \N__29516\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__5050\ : InMux
    port map (
            O => \N__29513\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__5049\ : InMux
    port map (
            O => \N__29510\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__5048\ : InMux
    port map (
            O => \N__29507\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__5047\ : InMux
    port map (
            O => \N__29504\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__5046\ : InMux
    port map (
            O => \N__29501\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__5045\ : InMux
    port map (
            O => \N__29498\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__5044\ : InMux
    port map (
            O => \N__29495\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__5043\ : InMux
    port map (
            O => \N__29492\,
            I => \bfn_11_12_0_\
        );

    \I__5042\ : InMux
    port map (
            O => \N__29489\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__5041\ : InMux
    port map (
            O => \N__29486\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__5040\ : InMux
    port map (
            O => \N__29483\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__5039\ : InMux
    port map (
            O => \N__29480\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__5038\ : InMux
    port map (
            O => \N__29477\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__5037\ : CascadeMux
    port map (
            O => \N__29474\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0_cascade_\
        );

    \I__5036\ : InMux
    port map (
            O => \N__29471\,
            I => \N__29465\
        );

    \I__5035\ : InMux
    port map (
            O => \N__29470\,
            I => \N__29465\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__29465\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__5033\ : InMux
    port map (
            O => \N__29462\,
            I => \N__29459\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__29459\,
            I => \N__29456\
        );

    \I__5031\ : Span4Mux_v
    port map (
            O => \N__29456\,
            I => \N__29450\
        );

    \I__5030\ : InMux
    port map (
            O => \N__29455\,
            I => \N__29443\
        );

    \I__5029\ : InMux
    port map (
            O => \N__29454\,
            I => \N__29443\
        );

    \I__5028\ : InMux
    port map (
            O => \N__29453\,
            I => \N__29443\
        );

    \I__5027\ : Odrv4
    port map (
            O => \N__29450\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__29443\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__5025\ : CascadeMux
    port map (
            O => \N__29438\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__5024\ : InMux
    port map (
            O => \N__29435\,
            I => \bfn_11_11_0_\
        );

    \I__5023\ : InMux
    port map (
            O => \N__29432\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__5022\ : InMux
    port map (
            O => \N__29429\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__5021\ : InMux
    port map (
            O => \N__29426\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__5020\ : InMux
    port map (
            O => \N__29423\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__5019\ : CascadeMux
    port map (
            O => \N__29420\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\
        );

    \I__5018\ : InMux
    port map (
            O => \N__29417\,
            I => \N__29413\
        );

    \I__5017\ : InMux
    port map (
            O => \N__29416\,
            I => \N__29409\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__29413\,
            I => \N__29406\
        );

    \I__5015\ : InMux
    port map (
            O => \N__29412\,
            I => \N__29403\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__29409\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__5013\ : Odrv4
    port map (
            O => \N__29406\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__29403\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__5011\ : InMux
    port map (
            O => \N__29396\,
            I => \N__29393\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__29393\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt16\
        );

    \I__5009\ : CascadeMux
    port map (
            O => \N__29390\,
            I => \N__29387\
        );

    \I__5008\ : InMux
    port map (
            O => \N__29387\,
            I => \N__29384\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__29384\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\
        );

    \I__5006\ : InMux
    port map (
            O => \N__29381\,
            I => \N__29378\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__29378\,
            I => \N__29375\
        );

    \I__5004\ : Span4Mux_h
    port map (
            O => \N__29375\,
            I => \N__29371\
        );

    \I__5003\ : InMux
    port map (
            O => \N__29374\,
            I => \N__29368\
        );

    \I__5002\ : Odrv4
    port map (
            O => \N__29371\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__29368\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__5000\ : CascadeMux
    port map (
            O => \N__29363\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17_cascade_\
        );

    \I__4999\ : CascadeMux
    port map (
            O => \N__29360\,
            I => \N__29357\
        );

    \I__4998\ : InMux
    port map (
            O => \N__29357\,
            I => \N__29351\
        );

    \I__4997\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29351\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__29351\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__4995\ : InMux
    port map (
            O => \N__29348\,
            I => \N__29345\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__29345\,
            I => \N__29341\
        );

    \I__4993\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29337\
        );

    \I__4992\ : Span4Mux_h
    port map (
            O => \N__29341\,
            I => \N__29334\
        );

    \I__4991\ : InMux
    port map (
            O => \N__29340\,
            I => \N__29331\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__29337\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__29334\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__29331\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__4987\ : InMux
    port map (
            O => \N__29324\,
            I => \N__29318\
        );

    \I__4986\ : InMux
    port map (
            O => \N__29323\,
            I => \N__29318\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__29318\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__4984\ : CascadeMux
    port map (
            O => \N__29315\,
            I => \N__29311\
        );

    \I__4983\ : InMux
    port map (
            O => \N__29314\,
            I => \N__29308\
        );

    \I__4982\ : InMux
    port map (
            O => \N__29311\,
            I => \N__29304\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__29308\,
            I => \N__29301\
        );

    \I__4980\ : InMux
    port map (
            O => \N__29307\,
            I => \N__29298\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__29304\,
            I => \N__29293\
        );

    \I__4978\ : Span4Mux_h
    port map (
            O => \N__29301\,
            I => \N__29293\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__29298\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__4976\ : Odrv4
    port map (
            O => \N__29293\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__4975\ : InMux
    port map (
            O => \N__29288\,
            I => \N__29285\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__29285\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__4973\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29279\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__29279\,
            I => \N__29276\
        );

    \I__4971\ : Odrv12
    port map (
            O => \N__29276\,
            I => \phase_controller_inst1.N_49_0\
        );

    \I__4970\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29267\
        );

    \I__4969\ : InMux
    port map (
            O => \N__29272\,
            I => \N__29264\
        );

    \I__4968\ : InMux
    port map (
            O => \N__29271\,
            I => \N__29259\
        );

    \I__4967\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29259\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__29267\,
            I => \N__29254\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__29264\,
            I => \N__29254\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__29259\,
            I => \N__29251\
        );

    \I__4963\ : Span4Mux_v
    port map (
            O => \N__29254\,
            I => \N__29248\
        );

    \I__4962\ : Span4Mux_h
    port map (
            O => \N__29251\,
            I => \N__29245\
        );

    \I__4961\ : Odrv4
    port map (
            O => \N__29248\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__4960\ : Odrv4
    port map (
            O => \N__29245\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__4959\ : InMux
    port map (
            O => \N__29240\,
            I => \N__29236\
        );

    \I__4958\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29233\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__29236\,
            I => \N__29230\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__29233\,
            I => \N__29225\
        );

    \I__4955\ : Span4Mux_v
    port map (
            O => \N__29230\,
            I => \N__29222\
        );

    \I__4954\ : InMux
    port map (
            O => \N__29229\,
            I => \N__29219\
        );

    \I__4953\ : InMux
    port map (
            O => \N__29228\,
            I => \N__29216\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__29225\,
            I => \N__29213\
        );

    \I__4951\ : Odrv4
    port map (
            O => \N__29222\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__29219\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__29216\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4948\ : Odrv4
    port map (
            O => \N__29213\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4947\ : InMux
    port map (
            O => \N__29204\,
            I => \N__29201\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__29201\,
            I => \N__29197\
        );

    \I__4945\ : InMux
    port map (
            O => \N__29200\,
            I => \N__29193\
        );

    \I__4944\ : Span4Mux_h
    port map (
            O => \N__29197\,
            I => \N__29190\
        );

    \I__4943\ : InMux
    port map (
            O => \N__29196\,
            I => \N__29187\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__29193\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__4941\ : Odrv4
    port map (
            O => \N__29190\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__29187\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__4939\ : InMux
    port map (
            O => \N__29180\,
            I => \N__29176\
        );

    \I__4938\ : InMux
    port map (
            O => \N__29179\,
            I => \N__29172\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__29176\,
            I => \N__29169\
        );

    \I__4936\ : InMux
    port map (
            O => \N__29175\,
            I => \N__29166\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__29172\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__4934\ : Odrv4
    port map (
            O => \N__29169\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__29166\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__4932\ : CascadeMux
    port map (
            O => \N__29159\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_\
        );

    \I__4931\ : InMux
    port map (
            O => \N__29156\,
            I => \N__29153\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__29153\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\
        );

    \I__4929\ : InMux
    port map (
            O => \N__29150\,
            I => \N__29147\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__29147\,
            I => \N__29144\
        );

    \I__4927\ : Odrv12
    port map (
            O => \N__29144\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\
        );

    \I__4926\ : InMux
    port map (
            O => \N__29141\,
            I => \N__29138\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__29138\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23\
        );

    \I__4924\ : CascadeMux
    port map (
            O => \N__29135\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_\
        );

    \I__4923\ : InMux
    port map (
            O => \N__29132\,
            I => \N__29129\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__29129\,
            I => \phase_controller_inst2.N_51_0\
        );

    \I__4921\ : InMux
    port map (
            O => \N__29126\,
            I => \N__29123\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__29123\,
            I => \N__29120\
        );

    \I__4919\ : Span4Mux_h
    port map (
            O => \N__29120\,
            I => \N__29114\
        );

    \I__4918\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29111\
        );

    \I__4917\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29108\
        );

    \I__4916\ : CascadeMux
    port map (
            O => \N__29117\,
            I => \N__29105\
        );

    \I__4915\ : Sp12to4
    port map (
            O => \N__29114\,
            I => \N__29098\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__29111\,
            I => \N__29098\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__29108\,
            I => \N__29098\
        );

    \I__4912\ : InMux
    port map (
            O => \N__29105\,
            I => \N__29095\
        );

    \I__4911\ : Span12Mux_v
    port map (
            O => \N__29098\,
            I => \N__29092\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__29095\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__4909\ : Odrv12
    port map (
            O => \N__29092\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__4908\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29080\
        );

    \I__4907\ : InMux
    port map (
            O => \N__29086\,
            I => \N__29080\
        );

    \I__4906\ : InMux
    port map (
            O => \N__29085\,
            I => \N__29077\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__29080\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__29077\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__29072\,
            I => \N__29069\
        );

    \I__4902\ : InMux
    port map (
            O => \N__29069\,
            I => \N__29065\
        );

    \I__4901\ : InMux
    port map (
            O => \N__29068\,
            I => \N__29062\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__29065\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__29062\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__4898\ : InMux
    port map (
            O => \N__29057\,
            I => \N__29054\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__29054\,
            I => \N__29051\
        );

    \I__4896\ : Odrv12
    port map (
            O => \N__29051\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__4895\ : InMux
    port map (
            O => \N__29048\,
            I => \N__29045\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__29045\,
            I => \N__29042\
        );

    \I__4893\ : Odrv12
    port map (
            O => \N__29042\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\
        );

    \I__4892\ : InMux
    port map (
            O => \N__29039\,
            I => \N__29036\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__29036\,
            I => \N__29033\
        );

    \I__4890\ : Odrv12
    port map (
            O => \N__29033\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\
        );

    \I__4889\ : InMux
    port map (
            O => \N__29030\,
            I => \N__29027\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__29027\,
            I => \N__29024\
        );

    \I__4887\ : Odrv12
    port map (
            O => \N__29024\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\
        );

    \I__4886\ : InMux
    port map (
            O => \N__29021\,
            I => \N__29016\
        );

    \I__4885\ : InMux
    port map (
            O => \N__29020\,
            I => \N__29012\
        );

    \I__4884\ : InMux
    port map (
            O => \N__29019\,
            I => \N__29009\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__29016\,
            I => \N__29006\
        );

    \I__4882\ : InMux
    port map (
            O => \N__29015\,
            I => \N__29003\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__29012\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__29009\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4879\ : Odrv12
    port map (
            O => \N__29006\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__29003\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4877\ : IoInMux
    port map (
            O => \N__28994\,
            I => \N__28991\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__28991\,
            I => \N__28988\
        );

    \I__4875\ : IoSpan4Mux
    port map (
            O => \N__28988\,
            I => \N__28985\
        );

    \I__4874\ : Span4Mux_s3_v
    port map (
            O => \N__28985\,
            I => \N__28982\
        );

    \I__4873\ : Span4Mux_v
    port map (
            O => \N__28982\,
            I => \N__28979\
        );

    \I__4872\ : Odrv4
    port map (
            O => \N__28979\,
            I => s4_phy_c
        );

    \I__4871\ : InMux
    port map (
            O => \N__28976\,
            I => \N__28971\
        );

    \I__4870\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28968\
        );

    \I__4869\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28965\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__28971\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__28968\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__28965\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__4865\ : InMux
    port map (
            O => \N__28958\,
            I => \N__28954\
        );

    \I__4864\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28950\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__28954\,
            I => \N__28947\
        );

    \I__4862\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28944\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__28950\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__4860\ : Odrv4
    port map (
            O => \N__28947\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__28944\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__4858\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28933\
        );

    \I__4857\ : InMux
    port map (
            O => \N__28936\,
            I => \N__28930\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__28933\,
            I => \N__28927\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__28930\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\
        );

    \I__4854\ : Odrv4
    port map (
            O => \N__28927\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\
        );

    \I__4853\ : CEMux
    port map (
            O => \N__28922\,
            I => \N__28889\
        );

    \I__4852\ : CEMux
    port map (
            O => \N__28921\,
            I => \N__28889\
        );

    \I__4851\ : CEMux
    port map (
            O => \N__28920\,
            I => \N__28889\
        );

    \I__4850\ : CEMux
    port map (
            O => \N__28919\,
            I => \N__28889\
        );

    \I__4849\ : CEMux
    port map (
            O => \N__28918\,
            I => \N__28889\
        );

    \I__4848\ : CEMux
    port map (
            O => \N__28917\,
            I => \N__28889\
        );

    \I__4847\ : CEMux
    port map (
            O => \N__28916\,
            I => \N__28889\
        );

    \I__4846\ : CEMux
    port map (
            O => \N__28915\,
            I => \N__28889\
        );

    \I__4845\ : CEMux
    port map (
            O => \N__28914\,
            I => \N__28889\
        );

    \I__4844\ : CEMux
    port map (
            O => \N__28913\,
            I => \N__28889\
        );

    \I__4843\ : CEMux
    port map (
            O => \N__28912\,
            I => \N__28889\
        );

    \I__4842\ : GlobalMux
    port map (
            O => \N__28889\,
            I => \N__28886\
        );

    \I__4841\ : gio2CtrlBuf
    port map (
            O => \N__28886\,
            I => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \I__4840\ : InMux
    port map (
            O => \N__28883\,
            I => \N__28878\
        );

    \I__4839\ : InMux
    port map (
            O => \N__28882\,
            I => \N__28873\
        );

    \I__4838\ : InMux
    port map (
            O => \N__28881\,
            I => \N__28873\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__28878\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__28873\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__4835\ : CascadeMux
    port map (
            O => \N__28868\,
            I => \N__28863\
        );

    \I__4834\ : InMux
    port map (
            O => \N__28867\,
            I => \N__28857\
        );

    \I__4833\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28857\
        );

    \I__4832\ : InMux
    port map (
            O => \N__28863\,
            I => \N__28852\
        );

    \I__4831\ : InMux
    port map (
            O => \N__28862\,
            I => \N__28852\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__28857\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__28852\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__4828\ : InMux
    port map (
            O => \N__28847\,
            I => \N__28844\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__28844\,
            I => \phase_controller_inst2.test_0_sqmuxa\
        );

    \I__4826\ : InMux
    port map (
            O => \N__28841\,
            I => \N__28838\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__28838\,
            I => \N__28835\
        );

    \I__4824\ : Span4Mux_v
    port map (
            O => \N__28835\,
            I => \N__28831\
        );

    \I__4823\ : InMux
    port map (
            O => \N__28834\,
            I => \N__28828\
        );

    \I__4822\ : Span4Mux_h
    port map (
            O => \N__28831\,
            I => \N__28825\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__28828\,
            I => \N__28822\
        );

    \I__4820\ : Span4Mux_v
    port map (
            O => \N__28825\,
            I => \N__28816\
        );

    \I__4819\ : Span4Mux_v
    port map (
            O => \N__28822\,
            I => \N__28813\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28808\
        );

    \I__4817\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28808\
        );

    \I__4816\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28805\
        );

    \I__4815\ : Span4Mux_v
    port map (
            O => \N__28816\,
            I => \N__28802\
        );

    \I__4814\ : Span4Mux_v
    port map (
            O => \N__28813\,
            I => \N__28795\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__28808\,
            I => \N__28795\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__28805\,
            I => \N__28795\
        );

    \I__4811\ : Odrv4
    port map (
            O => \N__28802\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__4810\ : Odrv4
    port map (
            O => \N__28795\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__4809\ : CascadeMux
    port map (
            O => \N__28790\,
            I => \N__28787\
        );

    \I__4808\ : InMux
    port map (
            O => \N__28787\,
            I => \N__28784\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__28784\,
            I => \N__28780\
        );

    \I__4806\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28777\
        );

    \I__4805\ : Span4Mux_v
    port map (
            O => \N__28780\,
            I => \N__28774\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__28777\,
            I => \N__28771\
        );

    \I__4803\ : Span4Mux_h
    port map (
            O => \N__28774\,
            I => \N__28768\
        );

    \I__4802\ : Span12Mux_s11_v
    port map (
            O => \N__28771\,
            I => \N__28763\
        );

    \I__4801\ : Span4Mux_v
    port map (
            O => \N__28768\,
            I => \N__28760\
        );

    \I__4800\ : InMux
    port map (
            O => \N__28767\,
            I => \N__28755\
        );

    \I__4799\ : InMux
    port map (
            O => \N__28766\,
            I => \N__28755\
        );

    \I__4798\ : Odrv12
    port map (
            O => \N__28763\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__28760\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__28755\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__4795\ : InMux
    port map (
            O => \N__28748\,
            I => \N__28744\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28747\,
            I => \N__28740\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__28744\,
            I => \N__28737\
        );

    \I__4792\ : InMux
    port map (
            O => \N__28743\,
            I => \N__28734\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__28740\,
            I => \N__28731\
        );

    \I__4790\ : Span4Mux_h
    port map (
            O => \N__28737\,
            I => \N__28728\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__28734\,
            I => \N__28725\
        );

    \I__4788\ : Span4Mux_v
    port map (
            O => \N__28731\,
            I => \N__28720\
        );

    \I__4787\ : Span4Mux_v
    port map (
            O => \N__28728\,
            I => \N__28720\
        );

    \I__4786\ : Span4Mux_h
    port map (
            O => \N__28725\,
            I => \N__28717\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__28720\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__4784\ : Odrv4
    port map (
            O => \N__28717\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__4783\ : InMux
    port map (
            O => \N__28712\,
            I => \N__28706\
        );

    \I__4782\ : InMux
    port map (
            O => \N__28711\,
            I => \N__28706\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__28706\,
            I => \N__28703\
        );

    \I__4780\ : Span4Mux_v
    port map (
            O => \N__28703\,
            I => \N__28699\
        );

    \I__4779\ : InMux
    port map (
            O => \N__28702\,
            I => \N__28696\
        );

    \I__4778\ : Span4Mux_h
    port map (
            O => \N__28699\,
            I => \N__28693\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__28696\,
            I => \N__28690\
        );

    \I__4776\ : Sp12to4
    port map (
            O => \N__28693\,
            I => \N__28685\
        );

    \I__4775\ : Span12Mux_h
    port map (
            O => \N__28690\,
            I => \N__28685\
        );

    \I__4774\ : Span12Mux_v
    port map (
            O => \N__28685\,
            I => \N__28682\
        );

    \I__4773\ : Odrv12
    port map (
            O => \N__28682\,
            I => il_min_comp2_c
        );

    \I__4772\ : InMux
    port map (
            O => \N__28679\,
            I => \N__28675\
        );

    \I__4771\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28672\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__28675\,
            I => \phase_controller_inst2.N_58\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__28672\,
            I => \phase_controller_inst2.N_58\
        );

    \I__4768\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28663\
        );

    \I__4767\ : InMux
    port map (
            O => \N__28666\,
            I => \N__28660\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__28663\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__28660\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__4764\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28651\
        );

    \I__4763\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28648\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__28651\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__28648\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__4760\ : InMux
    port map (
            O => \N__28643\,
            I => \N__28640\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__28640\,
            I => \N__28635\
        );

    \I__4758\ : InMux
    port map (
            O => \N__28639\,
            I => \N__28632\
        );

    \I__4757\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28629\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__28635\,
            I => \N__28626\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__28632\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__28629\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__28626\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4752\ : CascadeMux
    port map (
            O => \N__28619\,
            I => \N__28616\
        );

    \I__4751\ : InMux
    port map (
            O => \N__28616\,
            I => \N__28613\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__28613\,
            I => \N__28610\
        );

    \I__4749\ : Odrv12
    port map (
            O => \N__28610\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__4748\ : InMux
    port map (
            O => \N__28607\,
            I => \N__28604\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__28604\,
            I => \N__28601\
        );

    \I__4746\ : Odrv12
    port map (
            O => \N__28601\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__4745\ : InMux
    port map (
            O => \N__28598\,
            I => \N__28595\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__28595\,
            I => \N__28592\
        );

    \I__4743\ : Odrv12
    port map (
            O => \N__28592\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__4742\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28586\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__28586\,
            I => \N__28583\
        );

    \I__4740\ : Span4Mux_h
    port map (
            O => \N__28583\,
            I => \N__28579\
        );

    \I__4739\ : InMux
    port map (
            O => \N__28582\,
            I => \N__28575\
        );

    \I__4738\ : Sp12to4
    port map (
            O => \N__28579\,
            I => \N__28572\
        );

    \I__4737\ : InMux
    port map (
            O => \N__28578\,
            I => \N__28569\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__28575\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__4735\ : Odrv12
    port map (
            O => \N__28572\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__28569\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__4733\ : InMux
    port map (
            O => \N__28562\,
            I => \N__28557\
        );

    \I__4732\ : InMux
    port map (
            O => \N__28561\,
            I => \N__28554\
        );

    \I__4731\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28551\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__28557\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__28554\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__28551\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__4727\ : InMux
    port map (
            O => \N__28544\,
            I => \N__28538\
        );

    \I__4726\ : InMux
    port map (
            O => \N__28543\,
            I => \N__28538\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__28538\,
            I => \N__28535\
        );

    \I__4724\ : Span4Mux_v
    port map (
            O => \N__28535\,
            I => \N__28532\
        );

    \I__4723\ : Odrv4
    port map (
            O => \N__28532\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\
        );

    \I__4722\ : InMux
    port map (
            O => \N__28529\,
            I => \N__28523\
        );

    \I__4721\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28523\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__28523\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\
        );

    \I__4719\ : CascadeMux
    port map (
            O => \N__28520\,
            I => \N__28517\
        );

    \I__4718\ : InMux
    port map (
            O => \N__28517\,
            I => \N__28514\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__28514\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\
        );

    \I__4716\ : InMux
    port map (
            O => \N__28511\,
            I => \N__28508\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__28508\,
            I => \N__28503\
        );

    \I__4714\ : InMux
    port map (
            O => \N__28507\,
            I => \N__28500\
        );

    \I__4713\ : InMux
    port map (
            O => \N__28506\,
            I => \N__28497\
        );

    \I__4712\ : Span4Mux_v
    port map (
            O => \N__28503\,
            I => \N__28494\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__28500\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__28497\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__4709\ : Odrv4
    port map (
            O => \N__28494\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__4708\ : InMux
    port map (
            O => \N__28487\,
            I => \N__28484\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__28484\,
            I => \N__28481\
        );

    \I__4706\ : Odrv12
    port map (
            O => \N__28481\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__4705\ : InMux
    port map (
            O => \N__28478\,
            I => \N__28475\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__28475\,
            I => \N__28472\
        );

    \I__4703\ : Span4Mux_h
    port map (
            O => \N__28472\,
            I => \N__28468\
        );

    \I__4702\ : InMux
    port map (
            O => \N__28471\,
            I => \N__28465\
        );

    \I__4701\ : Odrv4
    port map (
            O => \N__28468\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__28465\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__4699\ : InMux
    port map (
            O => \N__28460\,
            I => \N__28457\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__28457\,
            I => \N__28454\
        );

    \I__4697\ : Span4Mux_v
    port map (
            O => \N__28454\,
            I => \N__28451\
        );

    \I__4696\ : Odrv4
    port map (
            O => \N__28451\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__28448\,
            I => \N__28445\
        );

    \I__4694\ : InMux
    port map (
            O => \N__28445\,
            I => \N__28442\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__28442\,
            I => \N__28439\
        );

    \I__4692\ : Odrv4
    port map (
            O => \N__28439\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt28\
        );

    \I__4691\ : InMux
    port map (
            O => \N__28436\,
            I => \N__28433\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__28433\,
            I => \N__28430\
        );

    \I__4689\ : Odrv4
    port map (
            O => \N__28430\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\
        );

    \I__4688\ : InMux
    port map (
            O => \N__28427\,
            I => \N__28424\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__28424\,
            I => \N__28421\
        );

    \I__4686\ : Span4Mux_h
    port map (
            O => \N__28421\,
            I => \N__28417\
        );

    \I__4685\ : InMux
    port map (
            O => \N__28420\,
            I => \N__28414\
        );

    \I__4684\ : Odrv4
    port map (
            O => \N__28417\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__28414\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__4682\ : CascadeMux
    port map (
            O => \N__28409\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29_cascade_\
        );

    \I__4681\ : CascadeMux
    port map (
            O => \N__28406\,
            I => \N__28403\
        );

    \I__4680\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28397\
        );

    \I__4679\ : InMux
    port map (
            O => \N__28402\,
            I => \N__28397\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__28397\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\
        );

    \I__4677\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28389\
        );

    \I__4676\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28386\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28383\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__28389\,
            I => \N__28380\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__28386\,
            I => \N__28377\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__28383\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__4671\ : Odrv12
    port map (
            O => \N__28380\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__4670\ : Odrv4
    port map (
            O => \N__28377\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__4669\ : InMux
    port map (
            O => \N__28370\,
            I => \N__28364\
        );

    \I__4668\ : InMux
    port map (
            O => \N__28369\,
            I => \N__28364\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__28364\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\
        );

    \I__4666\ : InMux
    port map (
            O => \N__28361\,
            I => \N__28358\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__28358\,
            I => \N__28355\
        );

    \I__4664\ : Odrv4
    port map (
            O => \N__28355\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt30\
        );

    \I__4663\ : InMux
    port map (
            O => \N__28352\,
            I => \N__28349\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__28349\,
            I => \N__28346\
        );

    \I__4661\ : Odrv12
    port map (
            O => \N__28346\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\
        );

    \I__4660\ : CascadeMux
    port map (
            O => \N__28343\,
            I => \N__28340\
        );

    \I__4659\ : InMux
    port map (
            O => \N__28340\,
            I => \N__28337\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__28337\,
            I => \N__28334\
        );

    \I__4657\ : Span4Mux_v
    port map (
            O => \N__28334\,
            I => \N__28331\
        );

    \I__4656\ : Odrv4
    port map (
            O => \N__28331\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt22\
        );

    \I__4655\ : InMux
    port map (
            O => \N__28328\,
            I => \N__28325\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__28325\,
            I => \N__28322\
        );

    \I__4653\ : Odrv4
    port map (
            O => \N__28322\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\
        );

    \I__4652\ : CascadeMux
    port map (
            O => \N__28319\,
            I => \N__28316\
        );

    \I__4651\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28313\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__28313\,
            I => \N__28310\
        );

    \I__4649\ : Odrv4
    port map (
            O => \N__28310\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt26\
        );

    \I__4648\ : CascadeMux
    port map (
            O => \N__28307\,
            I => \N__28304\
        );

    \I__4647\ : InMux
    port map (
            O => \N__28304\,
            I => \N__28301\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__28301\,
            I => \N__28298\
        );

    \I__4645\ : Span4Mux_h
    port map (
            O => \N__28298\,
            I => \N__28295\
        );

    \I__4644\ : Odrv4
    port map (
            O => \N__28295\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\
        );

    \I__4643\ : InMux
    port map (
            O => \N__28292\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30\
        );

    \I__4642\ : InMux
    port map (
            O => \N__28289\,
            I => \N__28286\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__28286\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt24\
        );

    \I__4640\ : CascadeMux
    port map (
            O => \N__28283\,
            I => \N__28280\
        );

    \I__4639\ : InMux
    port map (
            O => \N__28280\,
            I => \N__28277\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__28277\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__4637\ : InMux
    port map (
            O => \N__28274\,
            I => \N__28271\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__28271\,
            I => \N__28268\
        );

    \I__4635\ : Span4Mux_h
    port map (
            O => \N__28268\,
            I => \N__28265\
        );

    \I__4634\ : Odrv4
    port map (
            O => \N__28265\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__4633\ : CascadeMux
    port map (
            O => \N__28262\,
            I => \N__28259\
        );

    \I__4632\ : InMux
    port map (
            O => \N__28259\,
            I => \N__28256\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__28256\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__4630\ : InMux
    port map (
            O => \N__28253\,
            I => \N__28250\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__28250\,
            I => \N__28247\
        );

    \I__4628\ : Span4Mux_h
    port map (
            O => \N__28247\,
            I => \N__28244\
        );

    \I__4627\ : Odrv4
    port map (
            O => \N__28244\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__4626\ : CascadeMux
    port map (
            O => \N__28241\,
            I => \N__28238\
        );

    \I__4625\ : InMux
    port map (
            O => \N__28238\,
            I => \N__28235\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__28235\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__4623\ : CascadeMux
    port map (
            O => \N__28232\,
            I => \N__28229\
        );

    \I__4622\ : InMux
    port map (
            O => \N__28229\,
            I => \N__28226\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__28226\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__28223\,
            I => \N__28220\
        );

    \I__4619\ : InMux
    port map (
            O => \N__28220\,
            I => \N__28217\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__28217\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__28214\,
            I => \N__28211\
        );

    \I__4616\ : InMux
    port map (
            O => \N__28211\,
            I => \N__28208\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__28208\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__4614\ : InMux
    port map (
            O => \N__28205\,
            I => \N__28202\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__28202\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__4612\ : InMux
    port map (
            O => \N__28199\,
            I => \N__28196\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__28196\,
            I => \N__28193\
        );

    \I__4610\ : Odrv12
    port map (
            O => \N__28193\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__28190\,
            I => \N__28187\
        );

    \I__4608\ : InMux
    port map (
            O => \N__28187\,
            I => \N__28184\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__28184\,
            I => \N__28181\
        );

    \I__4606\ : Odrv12
    port map (
            O => \N__28181\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt18\
        );

    \I__4605\ : InMux
    port map (
            O => \N__28178\,
            I => \N__28175\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__28175\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt20\
        );

    \I__4603\ : CascadeMux
    port map (
            O => \N__28172\,
            I => \N__28169\
        );

    \I__4602\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28166\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__28166\,
            I => \N__28163\
        );

    \I__4600\ : Odrv4
    port map (
            O => \N__28163\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\
        );

    \I__4599\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28157\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__28157\,
            I => \N__28154\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__28154\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__4596\ : CascadeMux
    port map (
            O => \N__28151\,
            I => \N__28148\
        );

    \I__4595\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28145\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__28145\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__4593\ : InMux
    port map (
            O => \N__28142\,
            I => \N__28139\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__28139\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__28136\,
            I => \N__28133\
        );

    \I__4590\ : InMux
    port map (
            O => \N__28133\,
            I => \N__28130\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__28130\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__4588\ : InMux
    port map (
            O => \N__28127\,
            I => \N__28124\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__28124\,
            I => \N__28121\
        );

    \I__4586\ : Odrv4
    port map (
            O => \N__28121\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__4585\ : CascadeMux
    port map (
            O => \N__28118\,
            I => \N__28115\
        );

    \I__4584\ : InMux
    port map (
            O => \N__28115\,
            I => \N__28112\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__28112\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__4582\ : CascadeMux
    port map (
            O => \N__28109\,
            I => \N__28106\
        );

    \I__4581\ : InMux
    port map (
            O => \N__28106\,
            I => \N__28103\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__28103\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__4579\ : InMux
    port map (
            O => \N__28100\,
            I => \N__28097\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__28097\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__4577\ : CascadeMux
    port map (
            O => \N__28094\,
            I => \N__28091\
        );

    \I__4576\ : InMux
    port map (
            O => \N__28091\,
            I => \N__28088\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__28088\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__4574\ : CascadeMux
    port map (
            O => \N__28085\,
            I => \N__28082\
        );

    \I__4573\ : InMux
    port map (
            O => \N__28082\,
            I => \N__28079\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__28079\,
            I => \N__28076\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__28076\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__4570\ : InMux
    port map (
            O => \N__28073\,
            I => \N__28070\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__28070\,
            I => \N__28067\
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__28067\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__4567\ : CascadeMux
    port map (
            O => \N__28064\,
            I => \N__28061\
        );

    \I__4566\ : InMux
    port map (
            O => \N__28061\,
            I => \N__28058\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__28058\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__4564\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28052\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__28052\,
            I => \N__28049\
        );

    \I__4562\ : Odrv4
    port map (
            O => \N__28049\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__4561\ : InMux
    port map (
            O => \N__28046\,
            I => \N__28041\
        );

    \I__4560\ : InMux
    port map (
            O => \N__28045\,
            I => \N__28038\
        );

    \I__4559\ : InMux
    port map (
            O => \N__28044\,
            I => \N__28035\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__28041\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__28038\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__28035\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__4555\ : InMux
    port map (
            O => \N__28028\,
            I => \N__28023\
        );

    \I__4554\ : InMux
    port map (
            O => \N__28027\,
            I => \N__28020\
        );

    \I__4553\ : InMux
    port map (
            O => \N__28026\,
            I => \N__28017\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__28023\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__28020\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__28017\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__4549\ : InMux
    port map (
            O => \N__28010\,
            I => \N__28004\
        );

    \I__4548\ : InMux
    port map (
            O => \N__28009\,
            I => \N__28004\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__28004\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\
        );

    \I__4546\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27997\
        );

    \I__4545\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27994\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__27997\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__27994\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\
        );

    \I__4542\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27984\
        );

    \I__4541\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27981\
        );

    \I__4540\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27978\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__27984\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__27981\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__27978\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__4536\ : CascadeMux
    port map (
            O => \N__27971\,
            I => \N__27968\
        );

    \I__4535\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27965\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__27965\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__4533\ : InMux
    port map (
            O => \N__27962\,
            I => \N__27959\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__27959\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__4531\ : InMux
    port map (
            O => \N__27956\,
            I => \N__27953\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__27953\,
            I => \N__27950\
        );

    \I__4529\ : Odrv12
    port map (
            O => \N__27950\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\
        );

    \I__4528\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27944\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__27944\,
            I => \N__27941\
        );

    \I__4526\ : Odrv12
    port map (
            O => \N__27941\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__4525\ : IoInMux
    port map (
            O => \N__27938\,
            I => \N__27935\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__27935\,
            I => \N__27932\
        );

    \I__4523\ : Odrv12
    port map (
            O => \N__27932\,
            I => s3_phy_c
        );

    \I__4522\ : InMux
    port map (
            O => \N__27929\,
            I => \N__27926\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27923\
        );

    \I__4520\ : Glb2LocalMux
    port map (
            O => \N__27923\,
            I => \N__27920\
        );

    \I__4519\ : GlobalMux
    port map (
            O => \N__27920\,
            I => clk_12mhz
        );

    \I__4518\ : IoInMux
    port map (
            O => \N__27917\,
            I => \N__27914\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__27914\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__4516\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27905\
        );

    \I__4515\ : InMux
    port map (
            O => \N__27910\,
            I => \N__27905\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__27905\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__27902\,
            I => \N__27898\
        );

    \I__4512\ : InMux
    port map (
            O => \N__27901\,
            I => \N__27893\
        );

    \I__4511\ : InMux
    port map (
            O => \N__27898\,
            I => \N__27893\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__27893\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__4509\ : CascadeMux
    port map (
            O => \N__27890\,
            I => \N__27886\
        );

    \I__4508\ : InMux
    port map (
            O => \N__27889\,
            I => \N__27883\
        );

    \I__4507\ : InMux
    port map (
            O => \N__27886\,
            I => \N__27879\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__27883\,
            I => \N__27876\
        );

    \I__4505\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27873\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__27879\,
            I => \N__27870\
        );

    \I__4503\ : Span4Mux_h
    port map (
            O => \N__27876\,
            I => \N__27867\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__27873\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__4501\ : Odrv12
    port map (
            O => \N__27870\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__4500\ : Odrv4
    port map (
            O => \N__27867\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__4499\ : InMux
    port map (
            O => \N__27860\,
            I => \N__27855\
        );

    \I__4498\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27852\
        );

    \I__4497\ : InMux
    port map (
            O => \N__27858\,
            I => \N__27849\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__27855\,
            I => \N__27844\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__27852\,
            I => \N__27844\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__27849\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__27844\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__27839\,
            I => \N__27836\
        );

    \I__4491\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27833\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__27833\,
            I => \N__27830\
        );

    \I__4489\ : Odrv12
    port map (
            O => \N__27830\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__4488\ : InMux
    port map (
            O => \N__27827\,
            I => \N__27824\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__27824\,
            I => \N__27821\
        );

    \I__4486\ : Odrv12
    port map (
            O => \N__27821\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__4485\ : InMux
    port map (
            O => \N__27818\,
            I => \N__27815\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__27815\,
            I => \N__27812\
        );

    \I__4483\ : Odrv12
    port map (
            O => \N__27812\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\
        );

    \I__4482\ : CascadeMux
    port map (
            O => \N__27809\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__27806\,
            I => \N__27803\
        );

    \I__4480\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27797\
        );

    \I__4479\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27797\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__27797\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__4477\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27788\
        );

    \I__4476\ : InMux
    port map (
            O => \N__27793\,
            I => \N__27788\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27788\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\
        );

    \I__4474\ : InMux
    port map (
            O => \N__27785\,
            I => \N__27781\
        );

    \I__4473\ : InMux
    port map (
            O => \N__27784\,
            I => \N__27778\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__27781\,
            I => \N__27774\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__27778\,
            I => \N__27771\
        );

    \I__4470\ : InMux
    port map (
            O => \N__27777\,
            I => \N__27768\
        );

    \I__4469\ : Span4Mux_h
    port map (
            O => \N__27774\,
            I => \N__27763\
        );

    \I__4468\ : Span4Mux_v
    port map (
            O => \N__27771\,
            I => \N__27763\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__27768\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__27763\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__4465\ : CascadeMux
    port map (
            O => \N__27758\,
            I => \N__27754\
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__27757\,
            I => \N__27751\
        );

    \I__4463\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27748\
        );

    \I__4462\ : InMux
    port map (
            O => \N__27751\,
            I => \N__27745\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__27748\,
            I => \N__27741\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__27745\,
            I => \N__27738\
        );

    \I__4459\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27735\
        );

    \I__4458\ : Span4Mux_h
    port map (
            O => \N__27741\,
            I => \N__27732\
        );

    \I__4457\ : Span4Mux_v
    port map (
            O => \N__27738\,
            I => \N__27729\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__27735\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__4455\ : Odrv4
    port map (
            O => \N__27732\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__27729\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__27722\,
            I => \N__27719\
        );

    \I__4452\ : InMux
    port map (
            O => \N__27719\,
            I => \N__27716\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__27716\,
            I => \N__27713\
        );

    \I__4450\ : Odrv4
    port map (
            O => \N__27713\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt24\
        );

    \I__4449\ : InMux
    port map (
            O => \N__27710\,
            I => \N__27706\
        );

    \I__4448\ : InMux
    port map (
            O => \N__27709\,
            I => \N__27703\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__27706\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__27703\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\
        );

    \I__4445\ : InMux
    port map (
            O => \N__27698\,
            I => \N__27695\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__27695\,
            I => \N__27691\
        );

    \I__4443\ : InMux
    port map (
            O => \N__27694\,
            I => \N__27688\
        );

    \I__4442\ : Odrv4
    port map (
            O => \N__27691\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__27688\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\
        );

    \I__4440\ : InMux
    port map (
            O => \N__27683\,
            I => \N__27680\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__27680\,
            I => \N__27676\
        );

    \I__4438\ : InMux
    port map (
            O => \N__27679\,
            I => \N__27673\
        );

    \I__4437\ : Odrv12
    port map (
            O => \N__27676\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__27673\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\
        );

    \I__4435\ : InMux
    port map (
            O => \N__27668\,
            I => \N__27665\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__27665\,
            I => \N__27661\
        );

    \I__4433\ : InMux
    port map (
            O => \N__27664\,
            I => \N__27657\
        );

    \I__4432\ : Span4Mux_v
    port map (
            O => \N__27661\,
            I => \N__27654\
        );

    \I__4431\ : InMux
    port map (
            O => \N__27660\,
            I => \N__27651\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__27657\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4429\ : Odrv4
    port map (
            O => \N__27654\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__27651\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4427\ : InMux
    port map (
            O => \N__27644\,
            I => \N__27641\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__27641\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__4425\ : InMux
    port map (
            O => \N__27638\,
            I => \N__27635\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__27635\,
            I => \N__27631\
        );

    \I__4423\ : InMux
    port map (
            O => \N__27634\,
            I => \N__27628\
        );

    \I__4422\ : Odrv4
    port map (
            O => \N__27631\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__27628\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\
        );

    \I__4420\ : InMux
    port map (
            O => \N__27623\,
            I => \N__27619\
        );

    \I__4419\ : InMux
    port map (
            O => \N__27622\,
            I => \N__27616\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__27619\,
            I => \N__27613\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__27616\,
            I => \N__27610\
        );

    \I__4416\ : Span12Mux_v
    port map (
            O => \N__27613\,
            I => \N__27607\
        );

    \I__4415\ : Span4Mux_v
    port map (
            O => \N__27610\,
            I => \N__27604\
        );

    \I__4414\ : Odrv12
    port map (
            O => \N__27607\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\
        );

    \I__4413\ : Odrv4
    port map (
            O => \N__27604\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\
        );

    \I__4412\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27595\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__27598\,
            I => \N__27591\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__27595\,
            I => \N__27588\
        );

    \I__4409\ : InMux
    port map (
            O => \N__27594\,
            I => \N__27585\
        );

    \I__4408\ : InMux
    port map (
            O => \N__27591\,
            I => \N__27582\
        );

    \I__4407\ : Span4Mux_h
    port map (
            O => \N__27588\,
            I => \N__27579\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__27585\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__27582\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__4404\ : Odrv4
    port map (
            O => \N__27579\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__4403\ : CascadeMux
    port map (
            O => \N__27572\,
            I => \N__27569\
        );

    \I__4402\ : InMux
    port map (
            O => \N__27569\,
            I => \N__27566\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__27566\,
            I => \N__27561\
        );

    \I__4400\ : InMux
    port map (
            O => \N__27565\,
            I => \N__27558\
        );

    \I__4399\ : InMux
    port map (
            O => \N__27564\,
            I => \N__27555\
        );

    \I__4398\ : Span4Mux_h
    port map (
            O => \N__27561\,
            I => \N__27552\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__27558\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__27555\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__4395\ : Odrv4
    port map (
            O => \N__27552\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__4394\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27541\
        );

    \I__4393\ : InMux
    port map (
            O => \N__27544\,
            I => \N__27538\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__27541\,
            I => \N__27535\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__27538\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\
        );

    \I__4390\ : Odrv4
    port map (
            O => \N__27535\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\
        );

    \I__4389\ : InMux
    port map (
            O => \N__27530\,
            I => \N__27527\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__27527\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\
        );

    \I__4387\ : InMux
    port map (
            O => \N__27524\,
            I => \N__27521\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__27521\,
            I => \N__27516\
        );

    \I__4385\ : InMux
    port map (
            O => \N__27520\,
            I => \N__27513\
        );

    \I__4384\ : InMux
    port map (
            O => \N__27519\,
            I => \N__27510\
        );

    \I__4383\ : Span4Mux_h
    port map (
            O => \N__27516\,
            I => \N__27505\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__27513\,
            I => \N__27505\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__27510\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__27505\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__27500\,
            I => \N__27497\
        );

    \I__4378\ : InMux
    port map (
            O => \N__27497\,
            I => \N__27493\
        );

    \I__4377\ : CascadeMux
    port map (
            O => \N__27496\,
            I => \N__27490\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__27493\,
            I => \N__27486\
        );

    \I__4375\ : InMux
    port map (
            O => \N__27490\,
            I => \N__27483\
        );

    \I__4374\ : InMux
    port map (
            O => \N__27489\,
            I => \N__27480\
        );

    \I__4373\ : Span4Mux_h
    port map (
            O => \N__27486\,
            I => \N__27475\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__27483\,
            I => \N__27475\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__27480\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__4370\ : Odrv4
    port map (
            O => \N__27475\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__4369\ : InMux
    port map (
            O => \N__27470\,
            I => \N__27467\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__27467\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__4367\ : InMux
    port map (
            O => \N__27464\,
            I => \N__27460\
        );

    \I__4366\ : InMux
    port map (
            O => \N__27463\,
            I => \N__27457\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__27460\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__27457\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__4363\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27446\
        );

    \I__4362\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27446\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__27446\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__4360\ : CascadeMux
    port map (
            O => \N__27443\,
            I => \N__27440\
        );

    \I__4359\ : InMux
    port map (
            O => \N__27440\,
            I => \N__27434\
        );

    \I__4358\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27434\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__27434\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__27431\,
            I => \N__27428\
        );

    \I__4355\ : InMux
    port map (
            O => \N__27428\,
            I => \N__27425\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__27425\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__4353\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27419\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__27419\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__4351\ : InMux
    port map (
            O => \N__27416\,
            I => \N__27412\
        );

    \I__4350\ : InMux
    port map (
            O => \N__27415\,
            I => \N__27409\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__27412\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__27409\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__4347\ : CascadeMux
    port map (
            O => \N__27404\,
            I => \N__27401\
        );

    \I__4346\ : InMux
    port map (
            O => \N__27401\,
            I => \N__27398\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__27398\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__4344\ : InMux
    port map (
            O => \N__27395\,
            I => \N__27391\
        );

    \I__4343\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27387\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__27391\,
            I => \N__27384\
        );

    \I__4341\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27381\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__27387\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__27384\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__27381\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__4337\ : InMux
    port map (
            O => \N__27374\,
            I => \N__27371\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__27371\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__27368\,
            I => \N__27365\
        );

    \I__4334\ : InMux
    port map (
            O => \N__27365\,
            I => \N__27362\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__27362\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt22\
        );

    \I__4332\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27353\
        );

    \I__4331\ : InMux
    port map (
            O => \N__27358\,
            I => \N__27353\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__27353\,
            I => \N__27350\
        );

    \I__4329\ : Odrv12
    port map (
            O => \N__27350\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\
        );

    \I__4328\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27343\
        );

    \I__4327\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27340\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__27343\,
            I => \N__27335\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__27340\,
            I => \N__27335\
        );

    \I__4324\ : Odrv4
    port map (
            O => \N__27335\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\
        );

    \I__4323\ : CascadeMux
    port map (
            O => \N__27332\,
            I => \N__27329\
        );

    \I__4322\ : InMux
    port map (
            O => \N__27329\,
            I => \N__27325\
        );

    \I__4321\ : InMux
    port map (
            O => \N__27328\,
            I => \N__27322\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__27325\,
            I => \N__27316\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__27322\,
            I => \N__27316\
        );

    \I__4318\ : InMux
    port map (
            O => \N__27321\,
            I => \N__27313\
        );

    \I__4317\ : Span4Mux_h
    port map (
            O => \N__27316\,
            I => \N__27310\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__27313\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__4315\ : Odrv4
    port map (
            O => \N__27310\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__4314\ : CascadeMux
    port map (
            O => \N__27305\,
            I => \N__27301\
        );

    \I__4313\ : InMux
    port map (
            O => \N__27304\,
            I => \N__27296\
        );

    \I__4312\ : InMux
    port map (
            O => \N__27301\,
            I => \N__27296\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__27296\,
            I => \N__27292\
        );

    \I__4310\ : InMux
    port map (
            O => \N__27295\,
            I => \N__27289\
        );

    \I__4309\ : Span4Mux_h
    port map (
            O => \N__27292\,
            I => \N__27286\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__27289\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__4307\ : Odrv4
    port map (
            O => \N__27286\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__4306\ : InMux
    port map (
            O => \N__27281\,
            I => \N__27278\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__27278\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\
        );

    \I__4304\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27271\
        );

    \I__4303\ : InMux
    port map (
            O => \N__27274\,
            I => \N__27267\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__27271\,
            I => \N__27264\
        );

    \I__4301\ : InMux
    port map (
            O => \N__27270\,
            I => \N__27261\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__27267\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__4299\ : Odrv12
    port map (
            O => \N__27264\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__27261\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__4297\ : CascadeMux
    port map (
            O => \N__27254\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\
        );

    \I__4296\ : InMux
    port map (
            O => \N__27251\,
            I => \N__27248\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__27248\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt16\
        );

    \I__4294\ : InMux
    port map (
            O => \N__27245\,
            I => \N__27239\
        );

    \I__4293\ : InMux
    port map (
            O => \N__27244\,
            I => \N__27239\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__27239\,
            I => \N__27235\
        );

    \I__4291\ : InMux
    port map (
            O => \N__27238\,
            I => \N__27232\
        );

    \I__4290\ : Span4Mux_h
    port map (
            O => \N__27235\,
            I => \N__27229\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__27232\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__4288\ : Odrv4
    port map (
            O => \N__27229\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__4287\ : CascadeMux
    port map (
            O => \N__27224\,
            I => \N__27221\
        );

    \I__4286\ : InMux
    port map (
            O => \N__27221\,
            I => \N__27215\
        );

    \I__4285\ : InMux
    port map (
            O => \N__27220\,
            I => \N__27215\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__27215\,
            I => \N__27212\
        );

    \I__4283\ : Span4Mux_h
    port map (
            O => \N__27212\,
            I => \N__27208\
        );

    \I__4282\ : InMux
    port map (
            O => \N__27211\,
            I => \N__27205\
        );

    \I__4281\ : Span4Mux_h
    port map (
            O => \N__27208\,
            I => \N__27202\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__27205\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__4279\ : Odrv4
    port map (
            O => \N__27202\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__27197\,
            I => \N__27194\
        );

    \I__4277\ : InMux
    port map (
            O => \N__27194\,
            I => \N__27191\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__27191\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\
        );

    \I__4275\ : InMux
    port map (
            O => \N__27188\,
            I => \N__27184\
        );

    \I__4274\ : InMux
    port map (
            O => \N__27187\,
            I => \N__27181\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__27184\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__27181\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__4271\ : CascadeMux
    port map (
            O => \N__27176\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\
        );

    \I__4270\ : InMux
    port map (
            O => \N__27173\,
            I => \N__27169\
        );

    \I__4269\ : InMux
    port map (
            O => \N__27172\,
            I => \N__27166\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__27169\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__27166\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__27161\,
            I => \elapsed_time_ns_1_RNILK91B_0_9_cascade_\
        );

    \I__4265\ : InMux
    port map (
            O => \N__27158\,
            I => \N__27155\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__27155\,
            I => \N__27152\
        );

    \I__4263\ : Span4Mux_h
    port map (
            O => \N__27152\,
            I => \N__27149\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__27149\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\
        );

    \I__4261\ : InMux
    port map (
            O => \N__27146\,
            I => \N__27143\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__27143\,
            I => \N__27140\
        );

    \I__4259\ : Span4Mux_v
    port map (
            O => \N__27140\,
            I => \N__27137\
        );

    \I__4258\ : Span4Mux_h
    port map (
            O => \N__27137\,
            I => \N__27134\
        );

    \I__4257\ : Sp12to4
    port map (
            O => \N__27134\,
            I => \N__27131\
        );

    \I__4256\ : Span12Mux_h
    port map (
            O => \N__27131\,
            I => \N__27128\
        );

    \I__4255\ : Odrv12
    port map (
            O => \N__27128\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_15\
        );

    \I__4254\ : InMux
    port map (
            O => \N__27125\,
            I => \N__27122\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__27122\,
            I => \N__27117\
        );

    \I__4252\ : CascadeMux
    port map (
            O => \N__27121\,
            I => \N__27107\
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__27120\,
            I => \N__27104\
        );

    \I__4250\ : Span4Mux_v
    port map (
            O => \N__27117\,
            I => \N__27101\
        );

    \I__4249\ : CascadeMux
    port map (
            O => \N__27116\,
            I => \N__27098\
        );

    \I__4248\ : CascadeMux
    port map (
            O => \N__27115\,
            I => \N__27095\
        );

    \I__4247\ : CascadeMux
    port map (
            O => \N__27114\,
            I => \N__27091\
        );

    \I__4246\ : CascadeMux
    port map (
            O => \N__27113\,
            I => \N__27087\
        );

    \I__4245\ : CascadeMux
    port map (
            O => \N__27112\,
            I => \N__27084\
        );

    \I__4244\ : CascadeMux
    port map (
            O => \N__27111\,
            I => \N__27081\
        );

    \I__4243\ : CascadeMux
    port map (
            O => \N__27110\,
            I => \N__27078\
        );

    \I__4242\ : InMux
    port map (
            O => \N__27107\,
            I => \N__27073\
        );

    \I__4241\ : InMux
    port map (
            O => \N__27104\,
            I => \N__27073\
        );

    \I__4240\ : Span4Mux_h
    port map (
            O => \N__27101\,
            I => \N__27070\
        );

    \I__4239\ : InMux
    port map (
            O => \N__27098\,
            I => \N__27059\
        );

    \I__4238\ : InMux
    port map (
            O => \N__27095\,
            I => \N__27059\
        );

    \I__4237\ : InMux
    port map (
            O => \N__27094\,
            I => \N__27059\
        );

    \I__4236\ : InMux
    port map (
            O => \N__27091\,
            I => \N__27059\
        );

    \I__4235\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27059\
        );

    \I__4234\ : InMux
    port map (
            O => \N__27087\,
            I => \N__27054\
        );

    \I__4233\ : InMux
    port map (
            O => \N__27084\,
            I => \N__27054\
        );

    \I__4232\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27049\
        );

    \I__4231\ : InMux
    port map (
            O => \N__27078\,
            I => \N__27049\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__27073\,
            I => \N__27038\
        );

    \I__4229\ : Sp12to4
    port map (
            O => \N__27070\,
            I => \N__27038\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__27059\,
            I => \N__27038\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__27054\,
            I => \N__27038\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__27049\,
            I => \N__27038\
        );

    \I__4225\ : Span12Mux_v
    port map (
            O => \N__27038\,
            I => \N__27035\
        );

    \I__4224\ : Odrv12
    port map (
            O => \N__27035\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__4223\ : InMux
    port map (
            O => \N__27032\,
            I => \N__27029\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__27029\,
            I => \N__27026\
        );

    \I__4221\ : Span4Mux_h
    port map (
            O => \N__27026\,
            I => \N__27023\
        );

    \I__4220\ : Odrv4
    port map (
            O => \N__27023\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\
        );

    \I__4219\ : InMux
    port map (
            O => \N__27020\,
            I => \N__27017\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__27017\,
            I => \N__27014\
        );

    \I__4217\ : Odrv4
    port map (
            O => \N__27014\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__4216\ : InMux
    port map (
            O => \N__27011\,
            I => \N__27008\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__27008\,
            I => \N__27005\
        );

    \I__4214\ : Odrv12
    port map (
            O => \N__27005\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__4213\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26999\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__26999\,
            I => \N__26996\
        );

    \I__4211\ : Odrv4
    port map (
            O => \N__26996\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__4210\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26990\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__26990\,
            I => \N__26987\
        );

    \I__4208\ : Odrv4
    port map (
            O => \N__26987\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__4207\ : InMux
    port map (
            O => \N__26984\,
            I => \N__26981\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__26981\,
            I => \N__26978\
        );

    \I__4205\ : Odrv12
    port map (
            O => \N__26978\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\
        );

    \I__4204\ : CascadeMux
    port map (
            O => \N__26975\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8_cascade_\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__26972\,
            I => \N__26969\
        );

    \I__4202\ : InMux
    port map (
            O => \N__26969\,
            I => \N__26966\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__26966\,
            I => \N__26963\
        );

    \I__4200\ : Odrv12
    port map (
            O => \N__26963\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__4199\ : CascadeMux
    port map (
            O => \N__26960\,
            I => \N__26957\
        );

    \I__4198\ : InMux
    port map (
            O => \N__26957\,
            I => \N__26954\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__26954\,
            I => \N__26951\
        );

    \I__4196\ : Odrv4
    port map (
            O => \N__26951\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt26\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__26948\,
            I => \N__26943\
        );

    \I__4194\ : InMux
    port map (
            O => \N__26947\,
            I => \N__26940\
        );

    \I__4193\ : InMux
    port map (
            O => \N__26946\,
            I => \N__26935\
        );

    \I__4192\ : InMux
    port map (
            O => \N__26943\,
            I => \N__26935\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__26940\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__26935\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__4189\ : InMux
    port map (
            O => \N__26930\,
            I => \N__26925\
        );

    \I__4188\ : InMux
    port map (
            O => \N__26929\,
            I => \N__26920\
        );

    \I__4187\ : InMux
    port map (
            O => \N__26928\,
            I => \N__26920\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__26925\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__26920\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__4184\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26912\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__26912\,
            I => \N__26909\
        );

    \I__4182\ : Odrv4
    port map (
            O => \N__26909\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\
        );

    \I__4181\ : InMux
    port map (
            O => \N__26906\,
            I => \N__26900\
        );

    \I__4180\ : InMux
    port map (
            O => \N__26905\,
            I => \N__26900\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__26900\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__26897\,
            I => \N__26893\
        );

    \I__4177\ : InMux
    port map (
            O => \N__26896\,
            I => \N__26888\
        );

    \I__4176\ : InMux
    port map (
            O => \N__26893\,
            I => \N__26888\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__26888\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\
        );

    \I__4174\ : CascadeMux
    port map (
            O => \N__26885\,
            I => \N__26882\
        );

    \I__4173\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26879\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__26879\,
            I => \N__26876\
        );

    \I__4171\ : Span4Mux_h
    port map (
            O => \N__26876\,
            I => \N__26873\
        );

    \I__4170\ : Odrv4
    port map (
            O => \N__26873\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt28\
        );

    \I__4169\ : CascadeMux
    port map (
            O => \N__26870\,
            I => \N__26867\
        );

    \I__4168\ : InMux
    port map (
            O => \N__26867\,
            I => \N__26864\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__26864\,
            I => \N__26861\
        );

    \I__4166\ : Span4Mux_v
    port map (
            O => \N__26861\,
            I => \N__26858\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__26858\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26855\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30\
        );

    \I__4163\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26849\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__26849\,
            I => \N__26846\
        );

    \I__4161\ : Odrv4
    port map (
            O => \N__26846\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt20\
        );

    \I__4160\ : CascadeMux
    port map (
            O => \N__26843\,
            I => \N__26838\
        );

    \I__4159\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26835\
        );

    \I__4158\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26830\
        );

    \I__4157\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26830\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__26835\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__26830\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__4154\ : CascadeMux
    port map (
            O => \N__26825\,
            I => \N__26820\
        );

    \I__4153\ : InMux
    port map (
            O => \N__26824\,
            I => \N__26817\
        );

    \I__4152\ : InMux
    port map (
            O => \N__26823\,
            I => \N__26812\
        );

    \I__4151\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26812\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__26817\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__26812\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__26807\,
            I => \N__26804\
        );

    \I__4147\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26801\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__26801\,
            I => \N__26798\
        );

    \I__4145\ : Odrv4
    port map (
            O => \N__26798\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\
        );

    \I__4144\ : InMux
    port map (
            O => \N__26795\,
            I => \N__26789\
        );

    \I__4143\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26789\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__26789\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\
        );

    \I__4141\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26780\
        );

    \I__4140\ : InMux
    port map (
            O => \N__26785\,
            I => \N__26780\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__26780\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\
        );

    \I__4138\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26774\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__26774\,
            I => \N__26771\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__26771\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__4135\ : InMux
    port map (
            O => \N__26768\,
            I => \N__26764\
        );

    \I__4134\ : InMux
    port map (
            O => \N__26767\,
            I => \N__26761\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__26764\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__26761\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__4131\ : InMux
    port map (
            O => \N__26756\,
            I => \N__26753\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__26753\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__4129\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26746\
        );

    \I__4128\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26743\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__26746\,
            I => \N__26740\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__26743\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__26740\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__4124\ : CascadeMux
    port map (
            O => \N__26735\,
            I => \N__26732\
        );

    \I__4123\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26729\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__26729\,
            I => \N__26726\
        );

    \I__4121\ : Odrv4
    port map (
            O => \N__26726\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__4120\ : InMux
    port map (
            O => \N__26723\,
            I => \N__26719\
        );

    \I__4119\ : InMux
    port map (
            O => \N__26722\,
            I => \N__26716\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__26719\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__26716\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__4116\ : InMux
    port map (
            O => \N__26711\,
            I => \N__26708\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__26708\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__4114\ : InMux
    port map (
            O => \N__26705\,
            I => \N__26702\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__26702\,
            I => \N__26699\
        );

    \I__4112\ : Span4Mux_v
    port map (
            O => \N__26699\,
            I => \N__26696\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__26696\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__26693\,
            I => \N__26690\
        );

    \I__4109\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26687\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__26687\,
            I => \N__26684\
        );

    \I__4107\ : Span4Mux_v
    port map (
            O => \N__26684\,
            I => \N__26681\
        );

    \I__4106\ : Odrv4
    port map (
            O => \N__26681\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt18\
        );

    \I__4105\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26675\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__26675\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__4103\ : InMux
    port map (
            O => \N__26672\,
            I => \N__26668\
        );

    \I__4102\ : InMux
    port map (
            O => \N__26671\,
            I => \N__26665\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__26668\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__26665\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__4099\ : CascadeMux
    port map (
            O => \N__26660\,
            I => \N__26657\
        );

    \I__4098\ : InMux
    port map (
            O => \N__26657\,
            I => \N__26654\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__26654\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__4096\ : InMux
    port map (
            O => \N__26651\,
            I => \N__26647\
        );

    \I__4095\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26644\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__26647\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__26644\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__4092\ : CascadeMux
    port map (
            O => \N__26639\,
            I => \N__26636\
        );

    \I__4091\ : InMux
    port map (
            O => \N__26636\,
            I => \N__26633\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__26633\,
            I => \N__26630\
        );

    \I__4089\ : Odrv4
    port map (
            O => \N__26630\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__4088\ : InMux
    port map (
            O => \N__26627\,
            I => \N__26624\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__26624\,
            I => \N__26621\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__26621\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__4085\ : InMux
    port map (
            O => \N__26618\,
            I => \N__26614\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26617\,
            I => \N__26611\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__26614\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__26611\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__26606\,
            I => \N__26603\
        );

    \I__4080\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26600\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__26600\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__4078\ : InMux
    port map (
            O => \N__26597\,
            I => \N__26593\
        );

    \I__4077\ : InMux
    port map (
            O => \N__26596\,
            I => \N__26590\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__26593\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__26590\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__4074\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26582\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__26582\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__4072\ : InMux
    port map (
            O => \N__26579\,
            I => \N__26576\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__26576\,
            I => \N__26573\
        );

    \I__4070\ : Odrv4
    port map (
            O => \N__26573\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__4069\ : InMux
    port map (
            O => \N__26570\,
            I => \N__26566\
        );

    \I__4068\ : InMux
    port map (
            O => \N__26569\,
            I => \N__26563\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__26566\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__26563\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__4065\ : CascadeMux
    port map (
            O => \N__26558\,
            I => \N__26555\
        );

    \I__4064\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26552\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__26552\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__26549\,
            I => \N__26546\
        );

    \I__4061\ : InMux
    port map (
            O => \N__26546\,
            I => \N__26543\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__26543\,
            I => \N__26540\
        );

    \I__4059\ : Odrv12
    port map (
            O => \N__26540\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__4058\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26533\
        );

    \I__4057\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26530\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__26533\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__26530\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__4054\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26522\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__26522\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__4052\ : InMux
    port map (
            O => \N__26519\,
            I => \N__26515\
        );

    \I__4051\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26512\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__26515\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__26512\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__4048\ : InMux
    port map (
            O => \N__26507\,
            I => \N__26504\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__26504\,
            I => \N__26501\
        );

    \I__4046\ : Odrv12
    port map (
            O => \N__26501\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__26498\,
            I => \N__26495\
        );

    \I__4044\ : InMux
    port map (
            O => \N__26495\,
            I => \N__26492\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__26492\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__4042\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26485\
        );

    \I__4041\ : InMux
    port map (
            O => \N__26488\,
            I => \N__26482\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__26485\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__26482\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__4038\ : CascadeMux
    port map (
            O => \N__26477\,
            I => \N__26474\
        );

    \I__4037\ : InMux
    port map (
            O => \N__26474\,
            I => \N__26471\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__26471\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__4035\ : CascadeMux
    port map (
            O => \N__26468\,
            I => \N__26465\
        );

    \I__4034\ : InMux
    port map (
            O => \N__26465\,
            I => \N__26459\
        );

    \I__4033\ : InMux
    port map (
            O => \N__26464\,
            I => \N__26459\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__26459\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__4031\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26452\
        );

    \I__4030\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26449\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__26452\,
            I => \N__26444\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__26449\,
            I => \N__26444\
        );

    \I__4027\ : Span4Mux_h
    port map (
            O => \N__26444\,
            I => \N__26440\
        );

    \I__4026\ : CascadeMux
    port map (
            O => \N__26443\,
            I => \N__26437\
        );

    \I__4025\ : Span4Mux_v
    port map (
            O => \N__26440\,
            I => \N__26434\
        );

    \I__4024\ : InMux
    port map (
            O => \N__26437\,
            I => \N__26431\
        );

    \I__4023\ : Span4Mux_v
    port map (
            O => \N__26434\,
            I => \N__26428\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__26431\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__26428\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__26423\,
            I => \N__26420\
        );

    \I__4019\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26417\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__26417\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__4017\ : InMux
    port map (
            O => \N__26414\,
            I => \N__26410\
        );

    \I__4016\ : InMux
    port map (
            O => \N__26413\,
            I => \N__26407\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__26410\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__26407\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__4013\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26399\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__26399\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__4011\ : CascadeMux
    port map (
            O => \N__26396\,
            I => \N__26393\
        );

    \I__4010\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26390\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__26390\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__4008\ : InMux
    port map (
            O => \N__26387\,
            I => \N__26384\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__26384\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__4006\ : InMux
    port map (
            O => \N__26381\,
            I => \N__26377\
        );

    \I__4005\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26374\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__26377\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__26374\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__26369\,
            I => \N__26366\
        );

    \I__4001\ : InMux
    port map (
            O => \N__26366\,
            I => \N__26363\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__26363\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__26360\,
            I => \N__26357\
        );

    \I__3998\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26354\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__26354\,
            I => \N__26351\
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__26351\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__3995\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26344\
        );

    \I__3994\ : InMux
    port map (
            O => \N__26347\,
            I => \N__26341\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__26344\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__26341\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__3991\ : InMux
    port map (
            O => \N__26336\,
            I => \N__26333\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__26333\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__3989\ : InMux
    port map (
            O => \N__26330\,
            I => \N__26324\
        );

    \I__3988\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26324\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__26324\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__3986\ : InMux
    port map (
            O => \N__26321\,
            I => \N__26314\
        );

    \I__3985\ : InMux
    port map (
            O => \N__26320\,
            I => \N__26314\
        );

    \I__3984\ : InMux
    port map (
            O => \N__26319\,
            I => \N__26311\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__26314\,
            I => \N__26308\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__26311\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__3981\ : Odrv4
    port map (
            O => \N__26308\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__3980\ : CascadeMux
    port map (
            O => \N__26303\,
            I => \N__26300\
        );

    \I__3979\ : InMux
    port map (
            O => \N__26300\,
            I => \N__26293\
        );

    \I__3978\ : InMux
    port map (
            O => \N__26299\,
            I => \N__26293\
        );

    \I__3977\ : InMux
    port map (
            O => \N__26298\,
            I => \N__26290\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__26293\,
            I => \N__26287\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__26290\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__3974\ : Odrv4
    port map (
            O => \N__26287\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__3973\ : InMux
    port map (
            O => \N__26282\,
            I => \N__26279\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__26279\,
            I => \N__26276\
        );

    \I__3971\ : Odrv4
    port map (
            O => \N__26276\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__3970\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26270\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__26270\,
            I => \N__26267\
        );

    \I__3968\ : Odrv4
    port map (
            O => \N__26267\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__3967\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26261\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__26261\,
            I => \N__26258\
        );

    \I__3965\ : Odrv4
    port map (
            O => \N__26258\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__3964\ : InMux
    port map (
            O => \N__26255\,
            I => \N__26252\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__26252\,
            I => \N__26249\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__26249\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__3961\ : InMux
    port map (
            O => \N__26246\,
            I => \N__26243\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__26243\,
            I => \N__26240\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__26240\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__3958\ : InMux
    port map (
            O => \N__26237\,
            I => \N__26234\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__26234\,
            I => \N__26231\
        );

    \I__3956\ : Odrv12
    port map (
            O => \N__26231\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__3955\ : InMux
    port map (
            O => \N__26228\,
            I => \N__26225\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__26225\,
            I => \N__26222\
        );

    \I__3953\ : Span12Mux_v
    port map (
            O => \N__26222\,
            I => \N__26218\
        );

    \I__3952\ : InMux
    port map (
            O => \N__26221\,
            I => \N__26215\
        );

    \I__3951\ : Odrv12
    port map (
            O => \N__26218\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__26215\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__3949\ : IoInMux
    port map (
            O => \N__26210\,
            I => \N__26189\
        );

    \I__3948\ : InMux
    port map (
            O => \N__26209\,
            I => \N__26182\
        );

    \I__3947\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26182\
        );

    \I__3946\ : InMux
    port map (
            O => \N__26207\,
            I => \N__26182\
        );

    \I__3945\ : InMux
    port map (
            O => \N__26206\,
            I => \N__26162\
        );

    \I__3944\ : InMux
    port map (
            O => \N__26205\,
            I => \N__26162\
        );

    \I__3943\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26162\
        );

    \I__3942\ : InMux
    port map (
            O => \N__26203\,
            I => \N__26153\
        );

    \I__3941\ : InMux
    port map (
            O => \N__26202\,
            I => \N__26153\
        );

    \I__3940\ : InMux
    port map (
            O => \N__26201\,
            I => \N__26153\
        );

    \I__3939\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26153\
        );

    \I__3938\ : InMux
    port map (
            O => \N__26199\,
            I => \N__26144\
        );

    \I__3937\ : InMux
    port map (
            O => \N__26198\,
            I => \N__26144\
        );

    \I__3936\ : InMux
    port map (
            O => \N__26197\,
            I => \N__26144\
        );

    \I__3935\ : InMux
    port map (
            O => \N__26196\,
            I => \N__26144\
        );

    \I__3934\ : InMux
    port map (
            O => \N__26195\,
            I => \N__26135\
        );

    \I__3933\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26135\
        );

    \I__3932\ : InMux
    port map (
            O => \N__26193\,
            I => \N__26135\
        );

    \I__3931\ : InMux
    port map (
            O => \N__26192\,
            I => \N__26135\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__26189\,
            I => \N__26132\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__26182\,
            I => \N__26129\
        );

    \I__3928\ : InMux
    port map (
            O => \N__26181\,
            I => \N__26126\
        );

    \I__3927\ : InMux
    port map (
            O => \N__26180\,
            I => \N__26117\
        );

    \I__3926\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26117\
        );

    \I__3925\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26117\
        );

    \I__3924\ : InMux
    port map (
            O => \N__26177\,
            I => \N__26117\
        );

    \I__3923\ : InMux
    port map (
            O => \N__26176\,
            I => \N__26108\
        );

    \I__3922\ : InMux
    port map (
            O => \N__26175\,
            I => \N__26108\
        );

    \I__3921\ : InMux
    port map (
            O => \N__26174\,
            I => \N__26108\
        );

    \I__3920\ : InMux
    port map (
            O => \N__26173\,
            I => \N__26108\
        );

    \I__3919\ : InMux
    port map (
            O => \N__26172\,
            I => \N__26099\
        );

    \I__3918\ : InMux
    port map (
            O => \N__26171\,
            I => \N__26099\
        );

    \I__3917\ : InMux
    port map (
            O => \N__26170\,
            I => \N__26099\
        );

    \I__3916\ : InMux
    port map (
            O => \N__26169\,
            I => \N__26099\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__26162\,
            I => \N__26096\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__26153\,
            I => \N__26091\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__26144\,
            I => \N__26091\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__26135\,
            I => \N__26088\
        );

    \I__3911\ : Span12Mux_s2_v
    port map (
            O => \N__26132\,
            I => \N__26085\
        );

    \I__3910\ : Span12Mux_v
    port map (
            O => \N__26129\,
            I => \N__26080\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__26126\,
            I => \N__26080\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__26117\,
            I => \N__26067\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__26108\,
            I => \N__26067\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__26099\,
            I => \N__26067\
        );

    \I__3905\ : Span4Mux_v
    port map (
            O => \N__26096\,
            I => \N__26067\
        );

    \I__3904\ : Span4Mux_v
    port map (
            O => \N__26091\,
            I => \N__26067\
        );

    \I__3903\ : Span4Mux_h
    port map (
            O => \N__26088\,
            I => \N__26067\
        );

    \I__3902\ : Span12Mux_v
    port map (
            O => \N__26085\,
            I => \N__26064\
        );

    \I__3901\ : Odrv12
    port map (
            O => \N__26080\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__26067\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__3899\ : Odrv12
    port map (
            O => \N__26064\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__3898\ : InMux
    port map (
            O => \N__26057\,
            I => \N__26054\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__26054\,
            I => \N__26051\
        );

    \I__3896\ : Span4Mux_v
    port map (
            O => \N__26051\,
            I => \N__26048\
        );

    \I__3895\ : Odrv4
    port map (
            O => \N__26048\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__3894\ : InMux
    port map (
            O => \N__26045\,
            I => \N__26042\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__26042\,
            I => \N__26037\
        );

    \I__3892\ : InMux
    port map (
            O => \N__26041\,
            I => \N__26032\
        );

    \I__3891\ : InMux
    port map (
            O => \N__26040\,
            I => \N__26032\
        );

    \I__3890\ : Odrv12
    port map (
            O => \N__26037\,
            I => \current_shift_inst.PI_CTRL.N_160\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__26032\,
            I => \current_shift_inst.PI_CTRL.N_160\
        );

    \I__3888\ : InMux
    port map (
            O => \N__26027\,
            I => \N__26023\
        );

    \I__3887\ : InMux
    port map (
            O => \N__26026\,
            I => \N__26020\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__26023\,
            I => \N__26017\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__26020\,
            I => \N__26014\
        );

    \I__3884\ : Span4Mux_v
    port map (
            O => \N__26017\,
            I => \N__26009\
        );

    \I__3883\ : Span4Mux_s3_h
    port map (
            O => \N__26014\,
            I => \N__26009\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__26009\,
            I => \N__26006\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__26006\,
            I => pwm_duty_input_2
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__26003\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__26000\,
            I => \N__25997\
        );

    \I__3878\ : InMux
    port map (
            O => \N__25997\,
            I => \N__25992\
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__25996\,
            I => \N__25989\
        );

    \I__3876\ : InMux
    port map (
            O => \N__25995\,
            I => \N__25986\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__25992\,
            I => \N__25982\
        );

    \I__3874\ : InMux
    port map (
            O => \N__25989\,
            I => \N__25979\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__25986\,
            I => \N__25976\
        );

    \I__3872\ : InMux
    port map (
            O => \N__25985\,
            I => \N__25973\
        );

    \I__3871\ : Odrv12
    port map (
            O => \N__25982\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__25979\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__25976\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__25973\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3867\ : CascadeMux
    port map (
            O => \N__25964\,
            I => \N__25961\
        );

    \I__3866\ : InMux
    port map (
            O => \N__25961\,
            I => \N__25958\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__25958\,
            I => \N__25954\
        );

    \I__3864\ : InMux
    port map (
            O => \N__25957\,
            I => \N__25950\
        );

    \I__3863\ : Span4Mux_v
    port map (
            O => \N__25954\,
            I => \N__25946\
        );

    \I__3862\ : InMux
    port map (
            O => \N__25953\,
            I => \N__25943\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__25950\,
            I => \N__25940\
        );

    \I__3860\ : InMux
    port map (
            O => \N__25949\,
            I => \N__25937\
        );

    \I__3859\ : Odrv4
    port map (
            O => \N__25946\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__25943\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__3857\ : Odrv4
    port map (
            O => \N__25940\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__25937\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__25928\,
            I => \N__25925\
        );

    \I__3854\ : InMux
    port map (
            O => \N__25925\,
            I => \N__25921\
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__25924\,
            I => \N__25918\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__25921\,
            I => \N__25915\
        );

    \I__3851\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25911\
        );

    \I__3850\ : Span4Mux_v
    port map (
            O => \N__25915\,
            I => \N__25907\
        );

    \I__3849\ : InMux
    port map (
            O => \N__25914\,
            I => \N__25904\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__25911\,
            I => \N__25901\
        );

    \I__3847\ : InMux
    port map (
            O => \N__25910\,
            I => \N__25898\
        );

    \I__3846\ : Odrv4
    port map (
            O => \N__25907\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__25904\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3844\ : Odrv12
    port map (
            O => \N__25901\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__25898\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3842\ : CascadeMux
    port map (
            O => \N__25889\,
            I => \N__25886\
        );

    \I__3841\ : InMux
    port map (
            O => \N__25886\,
            I => \N__25883\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__25883\,
            I => \N__25878\
        );

    \I__3839\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25874\
        );

    \I__3838\ : CascadeMux
    port map (
            O => \N__25881\,
            I => \N__25871\
        );

    \I__3837\ : Span4Mux_v
    port map (
            O => \N__25878\,
            I => \N__25868\
        );

    \I__3836\ : InMux
    port map (
            O => \N__25877\,
            I => \N__25865\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__25874\,
            I => \N__25862\
        );

    \I__3834\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25859\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__25868\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__25865\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3831\ : Odrv4
    port map (
            O => \N__25862\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__25859\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__25850\,
            I => \N__25847\
        );

    \I__3828\ : InMux
    port map (
            O => \N__25847\,
            I => \N__25844\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__25844\,
            I => \N__25841\
        );

    \I__3826\ : Span4Mux_h
    port map (
            O => \N__25841\,
            I => \N__25838\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__25838\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25835\,
            I => \N__25832\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__25832\,
            I => \N__25829\
        );

    \I__3822\ : Span12Mux_s7_h
    port map (
            O => \N__25829\,
            I => \N__25826\
        );

    \I__3821\ : Odrv12
    port map (
            O => \N__25826\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__3820\ : InMux
    port map (
            O => \N__25823\,
            I => \N__25820\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__25820\,
            I => \N__25817\
        );

    \I__3818\ : Odrv4
    port map (
            O => \N__25817\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__3817\ : InMux
    port map (
            O => \N__25814\,
            I => \N__25811\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__25811\,
            I => \N__25808\
        );

    \I__3815\ : Span4Mux_h
    port map (
            O => \N__25808\,
            I => \N__25805\
        );

    \I__3814\ : Odrv4
    port map (
            O => \N__25805\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__3813\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25799\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__25799\,
            I => \N__25796\
        );

    \I__3811\ : Odrv12
    port map (
            O => \N__25796\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__3810\ : InMux
    port map (
            O => \N__25793\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__3809\ : InMux
    port map (
            O => \N__25790\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__3808\ : InMux
    port map (
            O => \N__25787\,
            I => \bfn_7_13_0_\
        );

    \I__3807\ : InMux
    port map (
            O => \N__25784\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__3806\ : InMux
    port map (
            O => \N__25781\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__3805\ : InMux
    port map (
            O => \N__25778\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__3804\ : InMux
    port map (
            O => \N__25775\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__3803\ : InMux
    port map (
            O => \N__25772\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__3802\ : InMux
    port map (
            O => \N__25769\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__3801\ : InMux
    port map (
            O => \N__25766\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__3800\ : InMux
    port map (
            O => \N__25763\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25760\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__3798\ : InMux
    port map (
            O => \N__25757\,
            I => \bfn_7_12_0_\
        );

    \I__3797\ : InMux
    port map (
            O => \N__25754\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__3796\ : InMux
    port map (
            O => \N__25751\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__3795\ : InMux
    port map (
            O => \N__25748\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__3794\ : InMux
    port map (
            O => \N__25745\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__3793\ : InMux
    port map (
            O => \N__25742\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__3792\ : InMux
    port map (
            O => \N__25739\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__3791\ : InMux
    port map (
            O => \N__25736\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__3790\ : InMux
    port map (
            O => \N__25733\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__3789\ : InMux
    port map (
            O => \N__25730\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__3788\ : InMux
    port map (
            O => \N__25727\,
            I => \bfn_7_11_0_\
        );

    \I__3787\ : InMux
    port map (
            O => \N__25724\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__3786\ : InMux
    port map (
            O => \N__25721\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__3785\ : InMux
    port map (
            O => \N__25718\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__3784\ : InMux
    port map (
            O => \N__25715\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__25712\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0_cascade_\
        );

    \I__3782\ : InMux
    port map (
            O => \N__25709\,
            I => \N__25703\
        );

    \I__3781\ : InMux
    port map (
            O => \N__25708\,
            I => \N__25703\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__25703\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__25700\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__25697\,
            I => \N__25694\
        );

    \I__3777\ : InMux
    port map (
            O => \N__25694\,
            I => \N__25691\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__25691\,
            I => \N__25688\
        );

    \I__3775\ : Odrv4
    port map (
            O => \N__25688\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\
        );

    \I__3774\ : InMux
    port map (
            O => \N__25685\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__3773\ : CascadeMux
    port map (
            O => \N__25682\,
            I => \N__25679\
        );

    \I__3772\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25676\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__25676\,
            I => \N__25673\
        );

    \I__3770\ : Odrv4
    port map (
            O => \N__25673\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30\
        );

    \I__3769\ : InMux
    port map (
            O => \N__25670\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__3768\ : InMux
    port map (
            O => \N__25667\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__3767\ : InMux
    port map (
            O => \N__25664\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__3766\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25657\
        );

    \I__3765\ : InMux
    port map (
            O => \N__25660\,
            I => \N__25654\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__25657\,
            I => \N__25651\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__25654\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__3762\ : Odrv4
    port map (
            O => \N__25651\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__3761\ : InMux
    port map (
            O => \N__25646\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__3760\ : InMux
    port map (
            O => \N__25643\,
            I => \N__25640\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__25640\,
            I => \N__25636\
        );

    \I__3758\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25633\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__25636\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__25633\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__3755\ : InMux
    port map (
            O => \N__25628\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__3754\ : CascadeMux
    port map (
            O => \N__25625\,
            I => \N__25622\
        );

    \I__3753\ : InMux
    port map (
            O => \N__25622\,
            I => \N__25619\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__25619\,
            I => \N__25613\
        );

    \I__3751\ : InMux
    port map (
            O => \N__25618\,
            I => \N__25610\
        );

    \I__3750\ : InMux
    port map (
            O => \N__25617\,
            I => \N__25607\
        );

    \I__3749\ : InMux
    port map (
            O => \N__25616\,
            I => \N__25604\
        );

    \I__3748\ : Span4Mux_v
    port map (
            O => \N__25613\,
            I => \N__25599\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__25610\,
            I => \N__25599\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__25607\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__25604\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__3744\ : Odrv4
    port map (
            O => \N__25599\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__3743\ : InMux
    port map (
            O => \N__25592\,
            I => \N__25589\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__25589\,
            I => \N__25585\
        );

    \I__3741\ : InMux
    port map (
            O => \N__25588\,
            I => \N__25582\
        );

    \I__3740\ : Odrv4
    port map (
            O => \N__25585\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__25582\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__3738\ : InMux
    port map (
            O => \N__25577\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__25574\,
            I => \N__25571\
        );

    \I__3736\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25568\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__25568\,
            I => \N__25564\
        );

    \I__3734\ : InMux
    port map (
            O => \N__25567\,
            I => \N__25560\
        );

    \I__3733\ : Span4Mux_v
    port map (
            O => \N__25564\,
            I => \N__25556\
        );

    \I__3732\ : InMux
    port map (
            O => \N__25563\,
            I => \N__25553\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__25560\,
            I => \N__25550\
        );

    \I__3730\ : InMux
    port map (
            O => \N__25559\,
            I => \N__25547\
        );

    \I__3729\ : Odrv4
    port map (
            O => \N__25556\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__25553\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__3727\ : Odrv4
    port map (
            O => \N__25550\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__25547\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__3725\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25534\
        );

    \I__3724\ : InMux
    port map (
            O => \N__25537\,
            I => \N__25531\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__25534\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__25531\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__3721\ : InMux
    port map (
            O => \N__25526\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__25523\,
            I => \N__25518\
        );

    \I__3719\ : InMux
    port map (
            O => \N__25522\,
            I => \N__25496\
        );

    \I__3718\ : InMux
    port map (
            O => \N__25521\,
            I => \N__25496\
        );

    \I__3717\ : InMux
    port map (
            O => \N__25518\,
            I => \N__25487\
        );

    \I__3716\ : InMux
    port map (
            O => \N__25517\,
            I => \N__25487\
        );

    \I__3715\ : InMux
    port map (
            O => \N__25516\,
            I => \N__25487\
        );

    \I__3714\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25487\
        );

    \I__3713\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25480\
        );

    \I__3712\ : InMux
    port map (
            O => \N__25513\,
            I => \N__25480\
        );

    \I__3711\ : InMux
    port map (
            O => \N__25512\,
            I => \N__25480\
        );

    \I__3710\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25476\
        );

    \I__3709\ : InMux
    port map (
            O => \N__25510\,
            I => \N__25467\
        );

    \I__3708\ : InMux
    port map (
            O => \N__25509\,
            I => \N__25462\
        );

    \I__3707\ : InMux
    port map (
            O => \N__25508\,
            I => \N__25462\
        );

    \I__3706\ : InMux
    port map (
            O => \N__25507\,
            I => \N__25447\
        );

    \I__3705\ : InMux
    port map (
            O => \N__25506\,
            I => \N__25447\
        );

    \I__3704\ : InMux
    port map (
            O => \N__25505\,
            I => \N__25447\
        );

    \I__3703\ : InMux
    port map (
            O => \N__25504\,
            I => \N__25447\
        );

    \I__3702\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25447\
        );

    \I__3701\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25447\
        );

    \I__3700\ : InMux
    port map (
            O => \N__25501\,
            I => \N__25447\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__25496\,
            I => \N__25440\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__25487\,
            I => \N__25440\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__25480\,
            I => \N__25440\
        );

    \I__3696\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25437\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__25476\,
            I => \N__25432\
        );

    \I__3694\ : InMux
    port map (
            O => \N__25475\,
            I => \N__25419\
        );

    \I__3693\ : InMux
    port map (
            O => \N__25474\,
            I => \N__25419\
        );

    \I__3692\ : InMux
    port map (
            O => \N__25473\,
            I => \N__25419\
        );

    \I__3691\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25419\
        );

    \I__3690\ : InMux
    port map (
            O => \N__25471\,
            I => \N__25419\
        );

    \I__3689\ : InMux
    port map (
            O => \N__25470\,
            I => \N__25419\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__25467\,
            I => \N__25414\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__25462\,
            I => \N__25414\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__25447\,
            I => \N__25409\
        );

    \I__3685\ : Span4Mux_v
    port map (
            O => \N__25440\,
            I => \N__25409\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__25437\,
            I => \N__25405\
        );

    \I__3683\ : InMux
    port map (
            O => \N__25436\,
            I => \N__25398\
        );

    \I__3682\ : InMux
    port map (
            O => \N__25435\,
            I => \N__25398\
        );

    \I__3681\ : Span12Mux_s10_v
    port map (
            O => \N__25432\,
            I => \N__25393\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__25419\,
            I => \N__25393\
        );

    \I__3679\ : Span4Mux_v
    port map (
            O => \N__25414\,
            I => \N__25390\
        );

    \I__3678\ : Sp12to4
    port map (
            O => \N__25409\,
            I => \N__25387\
        );

    \I__3677\ : InMux
    port map (
            O => \N__25408\,
            I => \N__25384\
        );

    \I__3676\ : Span4Mux_h
    port map (
            O => \N__25405\,
            I => \N__25381\
        );

    \I__3675\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25378\
        );

    \I__3674\ : InMux
    port map (
            O => \N__25403\,
            I => \N__25375\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__25398\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3672\ : Odrv12
    port map (
            O => \N__25393\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3671\ : Odrv4
    port map (
            O => \N__25390\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3670\ : Odrv12
    port map (
            O => \N__25387\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__25384\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__25381\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__25378\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__25375\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3665\ : InMux
    port map (
            O => \N__25358\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__25355\,
            I => \N__25350\
        );

    \I__3663\ : InMux
    port map (
            O => \N__25354\,
            I => \N__25347\
        );

    \I__3662\ : InMux
    port map (
            O => \N__25353\,
            I => \N__25344\
        );

    \I__3661\ : InMux
    port map (
            O => \N__25350\,
            I => \N__25341\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__25347\,
            I => \N__25338\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__25344\,
            I => \N__25335\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__25341\,
            I => \N__25332\
        );

    \I__3657\ : Span4Mux_h
    port map (
            O => \N__25338\,
            I => \N__25329\
        );

    \I__3656\ : Span4Mux_h
    port map (
            O => \N__25335\,
            I => \N__25326\
        );

    \I__3655\ : Odrv12
    port map (
            O => \N__25332\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__25329\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__25326\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__3652\ : InMux
    port map (
            O => \N__25319\,
            I => \N__25314\
        );

    \I__3651\ : InMux
    port map (
            O => \N__25318\,
            I => \N__25309\
        );

    \I__3650\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25309\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__25314\,
            I => \N__25306\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__25309\,
            I => \N__25303\
        );

    \I__3647\ : Span4Mux_s1_h
    port map (
            O => \N__25306\,
            I => \N__25300\
        );

    \I__3646\ : Span4Mux_v
    port map (
            O => \N__25303\,
            I => \N__25297\
        );

    \I__3645\ : Span4Mux_h
    port map (
            O => \N__25300\,
            I => \N__25294\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__25297\,
            I => pwm_duty_input_8
        );

    \I__3643\ : Odrv4
    port map (
            O => \N__25294\,
            I => pwm_duty_input_8
        );

    \I__3642\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25283\
        );

    \I__3641\ : InMux
    port map (
            O => \N__25288\,
            I => \N__25283\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__25283\,
            I => \N__25277\
        );

    \I__3639\ : InMux
    port map (
            O => \N__25282\,
            I => \N__25270\
        );

    \I__3638\ : InMux
    port map (
            O => \N__25281\,
            I => \N__25270\
        );

    \I__3637\ : InMux
    port map (
            O => \N__25280\,
            I => \N__25270\
        );

    \I__3636\ : Span4Mux_h
    port map (
            O => \N__25277\,
            I => \N__25263\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__25270\,
            I => \N__25263\
        );

    \I__3634\ : InMux
    port map (
            O => \N__25269\,
            I => \N__25260\
        );

    \I__3633\ : InMux
    port map (
            O => \N__25268\,
            I => \N__25257\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__25263\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__25260\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__25257\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__3629\ : InMux
    port map (
            O => \N__25250\,
            I => \N__25247\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__25247\,
            I => \N__25244\
        );

    \I__3627\ : Span4Mux_v
    port map (
            O => \N__25244\,
            I => \N__25237\
        );

    \I__3626\ : InMux
    port map (
            O => \N__25243\,
            I => \N__25228\
        );

    \I__3625\ : InMux
    port map (
            O => \N__25242\,
            I => \N__25228\
        );

    \I__3624\ : InMux
    port map (
            O => \N__25241\,
            I => \N__25228\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__25240\,
            I => \N__25224\
        );

    \I__3622\ : Span4Mux_v
    port map (
            O => \N__25237\,
            I => \N__25221\
        );

    \I__3621\ : InMux
    port map (
            O => \N__25236\,
            I => \N__25216\
        );

    \I__3620\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25216\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__25228\,
            I => \N__25211\
        );

    \I__3618\ : InMux
    port map (
            O => \N__25227\,
            I => \N__25206\
        );

    \I__3617\ : InMux
    port map (
            O => \N__25224\,
            I => \N__25206\
        );

    \I__3616\ : Span4Mux_v
    port map (
            O => \N__25221\,
            I => \N__25201\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__25216\,
            I => \N__25201\
        );

    \I__3614\ : InMux
    port map (
            O => \N__25215\,
            I => \N__25196\
        );

    \I__3613\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25196\
        );

    \I__3612\ : Span4Mux_v
    port map (
            O => \N__25211\,
            I => \N__25191\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__25206\,
            I => \N__25191\
        );

    \I__3610\ : Span4Mux_h
    port map (
            O => \N__25201\,
            I => \N__25188\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__25196\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__3608\ : Odrv4
    port map (
            O => \N__25191\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__25188\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__25181\,
            I => \N__25176\
        );

    \I__3605\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25171\
        );

    \I__3604\ : InMux
    port map (
            O => \N__25179\,
            I => \N__25171\
        );

    \I__3603\ : InMux
    port map (
            O => \N__25176\,
            I => \N__25168\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__25171\,
            I => \N__25165\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__25168\,
            I => \N__25162\
        );

    \I__3600\ : Span4Mux_h
    port map (
            O => \N__25165\,
            I => \N__25159\
        );

    \I__3599\ : Odrv12
    port map (
            O => \N__25162\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__25159\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__3597\ : CascadeMux
    port map (
            O => \N__25154\,
            I => \N__25148\
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__25153\,
            I => \N__25144\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__25152\,
            I => \N__25141\
        );

    \I__3594\ : InMux
    port map (
            O => \N__25151\,
            I => \N__25136\
        );

    \I__3593\ : InMux
    port map (
            O => \N__25148\,
            I => \N__25133\
        );

    \I__3592\ : InMux
    port map (
            O => \N__25147\,
            I => \N__25126\
        );

    \I__3591\ : InMux
    port map (
            O => \N__25144\,
            I => \N__25126\
        );

    \I__3590\ : InMux
    port map (
            O => \N__25141\,
            I => \N__25126\
        );

    \I__3589\ : InMux
    port map (
            O => \N__25140\,
            I => \N__25123\
        );

    \I__3588\ : InMux
    port map (
            O => \N__25139\,
            I => \N__25120\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__25136\,
            I => \current_shift_inst.PI_CTRL.N_158\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__25133\,
            I => \current_shift_inst.PI_CTRL.N_158\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__25126\,
            I => \current_shift_inst.PI_CTRL.N_158\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__25123\,
            I => \current_shift_inst.PI_CTRL.N_158\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__25120\,
            I => \current_shift_inst.PI_CTRL.N_158\
        );

    \I__3582\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25102\
        );

    \I__3581\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25102\
        );

    \I__3580\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25099\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__25102\,
            I => \N__25096\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__25099\,
            I => \N__25093\
        );

    \I__3577\ : Span4Mux_v
    port map (
            O => \N__25096\,
            I => \N__25090\
        );

    \I__3576\ : Span12Mux_s7_v
    port map (
            O => \N__25093\,
            I => \N__25087\
        );

    \I__3575\ : Odrv4
    port map (
            O => \N__25090\,
            I => pwm_duty_input_9
        );

    \I__3574\ : Odrv12
    port map (
            O => \N__25087\,
            I => pwm_duty_input_9
        );

    \I__3573\ : InMux
    port map (
            O => \N__25082\,
            I => \N__25079\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__25079\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__3570\ : InMux
    port map (
            O => \N__25073\,
            I => \N__25070\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__25070\,
            I => \N__25066\
        );

    \I__3568\ : CascadeMux
    port map (
            O => \N__25069\,
            I => \N__25061\
        );

    \I__3567\ : Span4Mux_v
    port map (
            O => \N__25066\,
            I => \N__25058\
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__25065\,
            I => \N__25055\
        );

    \I__3565\ : InMux
    port map (
            O => \N__25064\,
            I => \N__25052\
        );

    \I__3564\ : InMux
    port map (
            O => \N__25061\,
            I => \N__25049\
        );

    \I__3563\ : Span4Mux_v
    port map (
            O => \N__25058\,
            I => \N__25046\
        );

    \I__3562\ : InMux
    port map (
            O => \N__25055\,
            I => \N__25043\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__25052\,
            I => \N__25038\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__25049\,
            I => \N__25038\
        );

    \I__3559\ : Odrv4
    port map (
            O => \N__25046\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__25043\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__25038\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3556\ : InMux
    port map (
            O => \N__25031\,
            I => \N__25025\
        );

    \I__3555\ : InMux
    port map (
            O => \N__25030\,
            I => \N__25025\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__25025\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__3553\ : InMux
    port map (
            O => \N__25022\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__25019\,
            I => \N__25016\
        );

    \I__3551\ : InMux
    port map (
            O => \N__25016\,
            I => \N__25013\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__25013\,
            I => \N__25007\
        );

    \I__3549\ : InMux
    port map (
            O => \N__25012\,
            I => \N__25002\
        );

    \I__3548\ : InMux
    port map (
            O => \N__25011\,
            I => \N__25002\
        );

    \I__3547\ : InMux
    port map (
            O => \N__25010\,
            I => \N__24999\
        );

    \I__3546\ : Span12Mux_v
    port map (
            O => \N__25007\,
            I => \N__24994\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__25002\,
            I => \N__24994\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__24999\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3543\ : Odrv12
    port map (
            O => \N__24994\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__24989\,
            I => \N__24986\
        );

    \I__3541\ : InMux
    port map (
            O => \N__24986\,
            I => \N__24980\
        );

    \I__3540\ : InMux
    port map (
            O => \N__24985\,
            I => \N__24980\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__24980\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__3538\ : InMux
    port map (
            O => \N__24977\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__24974\,
            I => \N__24970\
        );

    \I__3536\ : CascadeMux
    port map (
            O => \N__24973\,
            I => \N__24967\
        );

    \I__3535\ : InMux
    port map (
            O => \N__24970\,
            I => \N__24964\
        );

    \I__3534\ : InMux
    port map (
            O => \N__24967\,
            I => \N__24959\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__24964\,
            I => \N__24956\
        );

    \I__3532\ : InMux
    port map (
            O => \N__24963\,
            I => \N__24953\
        );

    \I__3531\ : InMux
    port map (
            O => \N__24962\,
            I => \N__24950\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__24959\,
            I => \N__24943\
        );

    \I__3529\ : Sp12to4
    port map (
            O => \N__24956\,
            I => \N__24943\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__24953\,
            I => \N__24943\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__24950\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__3526\ : Odrv12
    port map (
            O => \N__24943\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__3525\ : InMux
    port map (
            O => \N__24938\,
            I => \N__24932\
        );

    \I__3524\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24932\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__24932\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__3522\ : InMux
    port map (
            O => \N__24929\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__24926\,
            I => \N__24923\
        );

    \I__3520\ : InMux
    port map (
            O => \N__24923\,
            I => \N__24920\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__24920\,
            I => \N__24917\
        );

    \I__3518\ : Span4Mux_h
    port map (
            O => \N__24917\,
            I => \N__24912\
        );

    \I__3517\ : InMux
    port map (
            O => \N__24916\,
            I => \N__24908\
        );

    \I__3516\ : InMux
    port map (
            O => \N__24915\,
            I => \N__24905\
        );

    \I__3515\ : Span4Mux_v
    port map (
            O => \N__24912\,
            I => \N__24902\
        );

    \I__3514\ : InMux
    port map (
            O => \N__24911\,
            I => \N__24899\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__24908\,
            I => \N__24894\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__24905\,
            I => \N__24894\
        );

    \I__3511\ : Odrv4
    port map (
            O => \N__24902\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__24899\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__24894\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3508\ : InMux
    port map (
            O => \N__24887\,
            I => \N__24881\
        );

    \I__3507\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24881\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__24881\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__3505\ : InMux
    port map (
            O => \N__24878\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__24875\,
            I => \N__24872\
        );

    \I__3503\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24869\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__24869\,
            I => \N__24866\
        );

    \I__3501\ : Span4Mux_h
    port map (
            O => \N__24866\,
            I => \N__24860\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__24865\,
            I => \N__24857\
        );

    \I__3499\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24854\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24863\,
            I => \N__24851\
        );

    \I__3497\ : Span4Mux_v
    port map (
            O => \N__24860\,
            I => \N__24848\
        );

    \I__3496\ : InMux
    port map (
            O => \N__24857\,
            I => \N__24845\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__24854\,
            I => \N__24840\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__24851\,
            I => \N__24840\
        );

    \I__3493\ : Odrv4
    port map (
            O => \N__24848\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__24845\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3491\ : Odrv4
    port map (
            O => \N__24840\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3490\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24827\
        );

    \I__3489\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24827\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__24827\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__3487\ : InMux
    port map (
            O => \N__24824\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__24821\,
            I => \N__24818\
        );

    \I__3485\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24815\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__24815\,
            I => \N__24811\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24814\,
            I => \N__24808\
        );

    \I__3482\ : Span4Mux_v
    port map (
            O => \N__24811\,
            I => \N__24803\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__24808\,
            I => \N__24800\
        );

    \I__3480\ : InMux
    port map (
            O => \N__24807\,
            I => \N__24795\
        );

    \I__3479\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24795\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__24803\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__24800\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__24795\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__24788\,
            I => \N__24784\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24787\,
            I => \N__24779\
        );

    \I__3473\ : InMux
    port map (
            O => \N__24784\,
            I => \N__24779\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__24779\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__3471\ : InMux
    port map (
            O => \N__24776\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\
        );

    \I__3470\ : InMux
    port map (
            O => \N__24773\,
            I => \N__24767\
        );

    \I__3469\ : InMux
    port map (
            O => \N__24772\,
            I => \N__24767\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__24767\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__3467\ : InMux
    port map (
            O => \N__24764\,
            I => \bfn_5_22_0_\
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__24761\,
            I => \N__24758\
        );

    \I__3465\ : InMux
    port map (
            O => \N__24758\,
            I => \N__24754\
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__24757\,
            I => \N__24751\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__24754\,
            I => \N__24748\
        );

    \I__3462\ : InMux
    port map (
            O => \N__24751\,
            I => \N__24745\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__24748\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__24745\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__24740\,
            I => \N__24737\
        );

    \I__3458\ : InMux
    port map (
            O => \N__24737\,
            I => \N__24734\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__24734\,
            I => \N__24730\
        );

    \I__3456\ : InMux
    port map (
            O => \N__24733\,
            I => \N__24727\
        );

    \I__3455\ : Span4Mux_h
    port map (
            O => \N__24730\,
            I => \N__24722\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__24727\,
            I => \N__24719\
        );

    \I__3453\ : InMux
    port map (
            O => \N__24726\,
            I => \N__24716\
        );

    \I__3452\ : InMux
    port map (
            O => \N__24725\,
            I => \N__24713\
        );

    \I__3451\ : Span4Mux_v
    port map (
            O => \N__24722\,
            I => \N__24710\
        );

    \I__3450\ : Span4Mux_v
    port map (
            O => \N__24719\,
            I => \N__24707\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__24716\,
            I => \N__24704\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__24713\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__3447\ : Odrv4
    port map (
            O => \N__24710\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__24707\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__3445\ : Odrv12
    port map (
            O => \N__24704\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__3444\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24689\
        );

    \I__3443\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24689\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__24689\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__3441\ : InMux
    port map (
            O => \N__24686\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__24683\,
            I => \N__24680\
        );

    \I__3439\ : InMux
    port map (
            O => \N__24680\,
            I => \N__24675\
        );

    \I__3438\ : InMux
    port map (
            O => \N__24679\,
            I => \N__24672\
        );

    \I__3437\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24669\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__24675\,
            I => \N__24663\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__24672\,
            I => \N__24663\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__24669\,
            I => \N__24660\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__24668\,
            I => \N__24657\
        );

    \I__3432\ : Span4Mux_v
    port map (
            O => \N__24663\,
            I => \N__24654\
        );

    \I__3431\ : Span4Mux_v
    port map (
            O => \N__24660\,
            I => \N__24651\
        );

    \I__3430\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24648\
        );

    \I__3429\ : Odrv4
    port map (
            O => \N__24654\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__24651\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__24648\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__3426\ : InMux
    port map (
            O => \N__24641\,
            I => \N__24635\
        );

    \I__3425\ : InMux
    port map (
            O => \N__24640\,
            I => \N__24635\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__24635\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__3423\ : InMux
    port map (
            O => \N__24632\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__24629\,
            I => \N__24624\
        );

    \I__3421\ : InMux
    port map (
            O => \N__24628\,
            I => \N__24621\
        );

    \I__3420\ : InMux
    port map (
            O => \N__24627\,
            I => \N__24618\
        );

    \I__3419\ : InMux
    port map (
            O => \N__24624\,
            I => \N__24615\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__24621\,
            I => \N__24609\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__24618\,
            I => \N__24609\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__24615\,
            I => \N__24606\
        );

    \I__3415\ : InMux
    port map (
            O => \N__24614\,
            I => \N__24603\
        );

    \I__3414\ : Span4Mux_v
    port map (
            O => \N__24609\,
            I => \N__24600\
        );

    \I__3413\ : Odrv12
    port map (
            O => \N__24606\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__24603\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__3411\ : Odrv4
    port map (
            O => \N__24600\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__24593\,
            I => \N__24589\
        );

    \I__3409\ : InMux
    port map (
            O => \N__24592\,
            I => \N__24586\
        );

    \I__3408\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24583\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__24586\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__24583\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__3405\ : InMux
    port map (
            O => \N__24578\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__24575\,
            I => \N__24572\
        );

    \I__3403\ : InMux
    port map (
            O => \N__24572\,
            I => \N__24568\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__24571\,
            I => \N__24565\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__24568\,
            I => \N__24561\
        );

    \I__3400\ : InMux
    port map (
            O => \N__24565\,
            I => \N__24558\
        );

    \I__3399\ : InMux
    port map (
            O => \N__24564\,
            I => \N__24555\
        );

    \I__3398\ : Span4Mux_v
    port map (
            O => \N__24561\,
            I => \N__24552\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__24558\,
            I => \N__24548\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__24555\,
            I => \N__24545\
        );

    \I__3395\ : Span4Mux_v
    port map (
            O => \N__24552\,
            I => \N__24542\
        );

    \I__3394\ : InMux
    port map (
            O => \N__24551\,
            I => \N__24539\
        );

    \I__3393\ : Span4Mux_s3_h
    port map (
            O => \N__24548\,
            I => \N__24534\
        );

    \I__3392\ : Span4Mux_v
    port map (
            O => \N__24545\,
            I => \N__24534\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__24542\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__24539\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__24534\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__3388\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24521\
        );

    \I__3387\ : InMux
    port map (
            O => \N__24526\,
            I => \N__24521\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__24521\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__3385\ : InMux
    port map (
            O => \N__24518\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__24515\,
            I => \N__24512\
        );

    \I__3383\ : InMux
    port map (
            O => \N__24512\,
            I => \N__24509\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__24509\,
            I => \N__24505\
        );

    \I__3381\ : CascadeMux
    port map (
            O => \N__24508\,
            I => \N__24502\
        );

    \I__3380\ : Span4Mux_h
    port map (
            O => \N__24505\,
            I => \N__24497\
        );

    \I__3379\ : InMux
    port map (
            O => \N__24502\,
            I => \N__24494\
        );

    \I__3378\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24491\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__24500\,
            I => \N__24488\
        );

    \I__3376\ : Span4Mux_h
    port map (
            O => \N__24497\,
            I => \N__24481\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__24494\,
            I => \N__24481\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__24491\,
            I => \N__24481\
        );

    \I__3373\ : InMux
    port map (
            O => \N__24488\,
            I => \N__24478\
        );

    \I__3372\ : Span4Mux_v
    port map (
            O => \N__24481\,
            I => \N__24475\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__24478\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3370\ : Odrv4
    port map (
            O => \N__24475\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3369\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24464\
        );

    \I__3368\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24464\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__24464\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__3366\ : InMux
    port map (
            O => \N__24461\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__3365\ : InMux
    port map (
            O => \N__24458\,
            I => \N__24455\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__24455\,
            I => \N__24450\
        );

    \I__3363\ : InMux
    port map (
            O => \N__24454\,
            I => \N__24447\
        );

    \I__3362\ : InMux
    port map (
            O => \N__24453\,
            I => \N__24443\
        );

    \I__3361\ : Span4Mux_v
    port map (
            O => \N__24450\,
            I => \N__24438\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__24447\,
            I => \N__24438\
        );

    \I__3359\ : InMux
    port map (
            O => \N__24446\,
            I => \N__24435\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__24443\,
            I => \N__24430\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__24438\,
            I => \N__24430\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__24435\,
            I => \N__24427\
        );

    \I__3355\ : Span4Mux_v
    port map (
            O => \N__24430\,
            I => \N__24424\
        );

    \I__3354\ : Odrv12
    port map (
            O => \N__24427\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__24424\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__24419\,
            I => \N__24415\
        );

    \I__3351\ : InMux
    port map (
            O => \N__24418\,
            I => \N__24410\
        );

    \I__3350\ : InMux
    port map (
            O => \N__24415\,
            I => \N__24410\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__24410\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__3348\ : InMux
    port map (
            O => \N__24407\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__24404\,
            I => \N__24401\
        );

    \I__3346\ : InMux
    port map (
            O => \N__24401\,
            I => \N__24397\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__24400\,
            I => \N__24393\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__24397\,
            I => \N__24389\
        );

    \I__3343\ : InMux
    port map (
            O => \N__24396\,
            I => \N__24386\
        );

    \I__3342\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24383\
        );

    \I__3341\ : InMux
    port map (
            O => \N__24392\,
            I => \N__24380\
        );

    \I__3340\ : Span4Mux_v
    port map (
            O => \N__24389\,
            I => \N__24377\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__24386\,
            I => \N__24374\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__24383\,
            I => \N__24369\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__24380\,
            I => \N__24369\
        );

    \I__3336\ : Odrv4
    port map (
            O => \N__24377\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3335\ : Odrv4
    port map (
            O => \N__24374\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3334\ : Odrv4
    port map (
            O => \N__24369\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__24362\,
            I => \N__24359\
        );

    \I__3332\ : InMux
    port map (
            O => \N__24359\,
            I => \N__24355\
        );

    \I__3331\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24352\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__24355\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__24352\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__3328\ : InMux
    port map (
            O => \N__24347\,
            I => \bfn_5_21_0_\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__24344\,
            I => \N__24341\
        );

    \I__3326\ : InMux
    port map (
            O => \N__24341\,
            I => \N__24338\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__24338\,
            I => \N__24334\
        );

    \I__3324\ : InMux
    port map (
            O => \N__24337\,
            I => \N__24330\
        );

    \I__3323\ : Span4Mux_h
    port map (
            O => \N__24334\,
            I => \N__24326\
        );

    \I__3322\ : InMux
    port map (
            O => \N__24333\,
            I => \N__24323\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__24330\,
            I => \N__24320\
        );

    \I__3320\ : InMux
    port map (
            O => \N__24329\,
            I => \N__24317\
        );

    \I__3319\ : Span4Mux_v
    port map (
            O => \N__24326\,
            I => \N__24310\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__24323\,
            I => \N__24310\
        );

    \I__3317\ : Span4Mux_v
    port map (
            O => \N__24320\,
            I => \N__24310\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__24317\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3315\ : Odrv4
    port map (
            O => \N__24310\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3314\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24301\
        );

    \I__3313\ : InMux
    port map (
            O => \N__24304\,
            I => \N__24298\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__24301\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__24298\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__3310\ : InMux
    port map (
            O => \N__24293\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__3309\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24287\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__24287\,
            I => \N__24284\
        );

    \I__3307\ : Odrv12
    port map (
            O => \N__24284\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__3306\ : CascadeMux
    port map (
            O => \N__24281\,
            I => \N__24278\
        );

    \I__3305\ : InMux
    port map (
            O => \N__24278\,
            I => \N__24273\
        );

    \I__3304\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24270\
        );

    \I__3303\ : InMux
    port map (
            O => \N__24276\,
            I => \N__24267\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__24273\,
            I => \N__24264\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__24270\,
            I => \N__24261\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__24267\,
            I => \N__24256\
        );

    \I__3299\ : Span4Mux_h
    port map (
            O => \N__24264\,
            I => \N__24256\
        );

    \I__3298\ : Span4Mux_v
    port map (
            O => \N__24261\,
            I => \N__24252\
        );

    \I__3297\ : Span4Mux_v
    port map (
            O => \N__24256\,
            I => \N__24249\
        );

    \I__3296\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24246\
        );

    \I__3295\ : Odrv4
    port map (
            O => \N__24252\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3294\ : Odrv4
    port map (
            O => \N__24249\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__24246\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3292\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24234\
        );

    \I__3291\ : InMux
    port map (
            O => \N__24238\,
            I => \N__24229\
        );

    \I__3290\ : InMux
    port map (
            O => \N__24237\,
            I => \N__24229\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__24234\,
            I => \N__24224\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__24229\,
            I => \N__24224\
        );

    \I__3287\ : Span4Mux_v
    port map (
            O => \N__24224\,
            I => \N__24221\
        );

    \I__3286\ : Odrv4
    port map (
            O => \N__24221\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__3285\ : InMux
    port map (
            O => \N__24218\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__3284\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24212\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__24212\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__24209\,
            I => \N__24204\
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__24208\,
            I => \N__24201\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__24207\,
            I => \N__24198\
        );

    \I__3279\ : InMux
    port map (
            O => \N__24204\,
            I => \N__24194\
        );

    \I__3278\ : InMux
    port map (
            O => \N__24201\,
            I => \N__24191\
        );

    \I__3277\ : InMux
    port map (
            O => \N__24198\,
            I => \N__24188\
        );

    \I__3276\ : InMux
    port map (
            O => \N__24197\,
            I => \N__24185\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__24194\,
            I => \N__24182\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__24191\,
            I => \N__24179\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__24188\,
            I => \N__24176\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__24185\,
            I => \N__24173\
        );

    \I__3271\ : Span4Mux_v
    port map (
            O => \N__24182\,
            I => \N__24170\
        );

    \I__3270\ : Span4Mux_h
    port map (
            O => \N__24179\,
            I => \N__24167\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__24176\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__24173\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3267\ : Odrv4
    port map (
            O => \N__24170\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3266\ : Odrv4
    port map (
            O => \N__24167\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3265\ : InMux
    port map (
            O => \N__24158\,
            I => \N__24152\
        );

    \I__3264\ : InMux
    port map (
            O => \N__24157\,
            I => \N__24149\
        );

    \I__3263\ : InMux
    port map (
            O => \N__24156\,
            I => \N__24144\
        );

    \I__3262\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24144\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__24152\,
            I => \N__24139\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__24149\,
            I => \N__24139\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__24144\,
            I => \N__24136\
        );

    \I__3258\ : Span4Mux_v
    port map (
            O => \N__24139\,
            I => \N__24133\
        );

    \I__3257\ : Span4Mux_h
    port map (
            O => \N__24136\,
            I => \N__24130\
        );

    \I__3256\ : Odrv4
    port map (
            O => \N__24133\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__3255\ : Odrv4
    port map (
            O => \N__24130\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__3254\ : InMux
    port map (
            O => \N__24125\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__3253\ : InMux
    port map (
            O => \N__24122\,
            I => \N__24119\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__24119\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__24116\,
            I => \N__24112\
        );

    \I__3250\ : InMux
    port map (
            O => \N__24115\,
            I => \N__24108\
        );

    \I__3249\ : InMux
    port map (
            O => \N__24112\,
            I => \N__24105\
        );

    \I__3248\ : InMux
    port map (
            O => \N__24111\,
            I => \N__24101\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__24108\,
            I => \N__24098\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__24105\,
            I => \N__24095\
        );

    \I__3245\ : InMux
    port map (
            O => \N__24104\,
            I => \N__24092\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__24101\,
            I => \N__24089\
        );

    \I__3243\ : Span4Mux_v
    port map (
            O => \N__24098\,
            I => \N__24086\
        );

    \I__3242\ : Span12Mux_h
    port map (
            O => \N__24095\,
            I => \N__24081\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__24092\,
            I => \N__24081\
        );

    \I__3240\ : Span4Mux_h
    port map (
            O => \N__24089\,
            I => \N__24078\
        );

    \I__3239\ : Odrv4
    port map (
            O => \N__24086\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3238\ : Odrv12
    port map (
            O => \N__24081\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__24078\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__24071\,
            I => \N__24067\
        );

    \I__3235\ : InMux
    port map (
            O => \N__24070\,
            I => \N__24063\
        );

    \I__3234\ : InMux
    port map (
            O => \N__24067\,
            I => \N__24060\
        );

    \I__3233\ : InMux
    port map (
            O => \N__24066\,
            I => \N__24057\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__24063\,
            I => \N__24054\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__24060\,
            I => \N__24051\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__24057\,
            I => \N__24048\
        );

    \I__3229\ : Span4Mux_v
    port map (
            O => \N__24054\,
            I => \N__24045\
        );

    \I__3228\ : Span4Mux_h
    port map (
            O => \N__24051\,
            I => \N__24042\
        );

    \I__3227\ : Span4Mux_h
    port map (
            O => \N__24048\,
            I => \N__24039\
        );

    \I__3226\ : Odrv4
    port map (
            O => \N__24045\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__3225\ : Odrv4
    port map (
            O => \N__24042\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__3224\ : Odrv4
    port map (
            O => \N__24039\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__3223\ : InMux
    port map (
            O => \N__24032\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__3222\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24025\
        );

    \I__3221\ : CascadeMux
    port map (
            O => \N__24028\,
            I => \N__24021\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__24025\,
            I => \N__24018\
        );

    \I__3219\ : InMux
    port map (
            O => \N__24024\,
            I => \N__24015\
        );

    \I__3218\ : InMux
    port map (
            O => \N__24021\,
            I => \N__24012\
        );

    \I__3217\ : Span4Mux_v
    port map (
            O => \N__24018\,
            I => \N__24007\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__24015\,
            I => \N__24007\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__24012\,
            I => \N__24004\
        );

    \I__3214\ : Span4Mux_v
    port map (
            O => \N__24007\,
            I => \N__23998\
        );

    \I__3213\ : Span4Mux_h
    port map (
            O => \N__24004\,
            I => \N__23998\
        );

    \I__3212\ : InMux
    port map (
            O => \N__24003\,
            I => \N__23995\
        );

    \I__3211\ : Span4Mux_v
    port map (
            O => \N__23998\,
            I => \N__23992\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__23995\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__23992\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__23987\,
            I => \N__23984\
        );

    \I__3207\ : InMux
    port map (
            O => \N__23984\,
            I => \N__23981\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__23981\,
            I => \N__23978\
        );

    \I__3205\ : Odrv4
    port map (
            O => \N__23978\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__3204\ : InMux
    port map (
            O => \N__23975\,
            I => \N__23970\
        );

    \I__3203\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23965\
        );

    \I__3202\ : InMux
    port map (
            O => \N__23973\,
            I => \N__23965\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__23970\,
            I => \N__23962\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__23965\,
            I => \N__23959\
        );

    \I__3199\ : Span4Mux_v
    port map (
            O => \N__23962\,
            I => \N__23956\
        );

    \I__3198\ : Span4Mux_h
    port map (
            O => \N__23959\,
            I => \N__23953\
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__23956\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__3196\ : Odrv4
    port map (
            O => \N__23953\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__3195\ : InMux
    port map (
            O => \N__23948\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__3194\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23942\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__23942\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__23939\,
            I => \N__23936\
        );

    \I__3191\ : InMux
    port map (
            O => \N__23936\,
            I => \N__23933\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__23933\,
            I => \N__23928\
        );

    \I__3189\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23925\
        );

    \I__3188\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23922\
        );

    \I__3187\ : Span4Mux_h
    port map (
            O => \N__23928\,
            I => \N__23914\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__23925\,
            I => \N__23914\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__23922\,
            I => \N__23914\
        );

    \I__3184\ : InMux
    port map (
            O => \N__23921\,
            I => \N__23911\
        );

    \I__3183\ : Span4Mux_v
    port map (
            O => \N__23914\,
            I => \N__23908\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__23911\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3181\ : Odrv4
    port map (
            O => \N__23908\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3180\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23898\
        );

    \I__3179\ : InMux
    port map (
            O => \N__23902\,
            I => \N__23895\
        );

    \I__3178\ : InMux
    port map (
            O => \N__23901\,
            I => \N__23892\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__23898\,
            I => \N__23889\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__23895\,
            I => \N__23886\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__23892\,
            I => \N__23883\
        );

    \I__3174\ : Span4Mux_v
    port map (
            O => \N__23889\,
            I => \N__23880\
        );

    \I__3173\ : Span4Mux_h
    port map (
            O => \N__23886\,
            I => \N__23877\
        );

    \I__3172\ : Span4Mux_h
    port map (
            O => \N__23883\,
            I => \N__23874\
        );

    \I__3171\ : Odrv4
    port map (
            O => \N__23880\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__3170\ : Odrv4
    port map (
            O => \N__23877\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__3169\ : Odrv4
    port map (
            O => \N__23874\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__3168\ : InMux
    port map (
            O => \N__23867\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__3167\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23861\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__23861\,
            I => \N__23858\
        );

    \I__3165\ : Odrv4
    port map (
            O => \N__23858\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__23855\,
            I => \N__23852\
        );

    \I__3163\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23849\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__23849\,
            I => \N__23844\
        );

    \I__3161\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23841\
        );

    \I__3160\ : InMux
    port map (
            O => \N__23847\,
            I => \N__23838\
        );

    \I__3159\ : Span4Mux_v
    port map (
            O => \N__23844\,
            I => \N__23835\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__23841\,
            I => \N__23829\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__23838\,
            I => \N__23829\
        );

    \I__3156\ : Span4Mux_v
    port map (
            O => \N__23835\,
            I => \N__23826\
        );

    \I__3155\ : InMux
    port map (
            O => \N__23834\,
            I => \N__23823\
        );

    \I__3154\ : Span4Mux_v
    port map (
            O => \N__23829\,
            I => \N__23820\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__23826\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__23823\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3151\ : Odrv4
    port map (
            O => \N__23820\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23813\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\
        );

    \I__3149\ : CascadeMux
    port map (
            O => \N__23810\,
            I => \N__23807\
        );

    \I__3148\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23803\
        );

    \I__3147\ : InMux
    port map (
            O => \N__23806\,
            I => \N__23800\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__23803\,
            I => \N__23797\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__23800\,
            I => \N__23793\
        );

    \I__3144\ : Span4Mux_h
    port map (
            O => \N__23797\,
            I => \N__23790\
        );

    \I__3143\ : InMux
    port map (
            O => \N__23796\,
            I => \N__23786\
        );

    \I__3142\ : Span4Mux_v
    port map (
            O => \N__23793\,
            I => \N__23783\
        );

    \I__3141\ : Span4Mux_v
    port map (
            O => \N__23790\,
            I => \N__23780\
        );

    \I__3140\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23777\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__23786\,
            I => \N__23774\
        );

    \I__3138\ : Odrv4
    port map (
            O => \N__23783\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3137\ : Odrv4
    port map (
            O => \N__23780\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__23777\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3135\ : Odrv12
    port map (
            O => \N__23774\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23765\,
            I => \bfn_5_20_0_\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__23762\,
            I => \N__23758\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__23761\,
            I => \N__23754\
        );

    \I__3131\ : InMux
    port map (
            O => \N__23758\,
            I => \N__23751\
        );

    \I__3130\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23748\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23754\,
            I => \N__23745\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__23751\,
            I => \N__23742\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__23748\,
            I => \N__23737\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__23745\,
            I => \N__23737\
        );

    \I__3125\ : Span4Mux_v
    port map (
            O => \N__23742\,
            I => \N__23731\
        );

    \I__3124\ : Span4Mux_v
    port map (
            O => \N__23737\,
            I => \N__23731\
        );

    \I__3123\ : InMux
    port map (
            O => \N__23736\,
            I => \N__23728\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__23731\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__23728\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3120\ : InMux
    port map (
            O => \N__23723\,
            I => \N__23717\
        );

    \I__3119\ : InMux
    port map (
            O => \N__23722\,
            I => \N__23717\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__23717\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__3117\ : InMux
    port map (
            O => \N__23714\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__23711\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\
        );

    \I__3115\ : InMux
    port map (
            O => \N__23708\,
            I => \N__23705\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__23705\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__3113\ : InMux
    port map (
            O => \N__23702\,
            I => \N__23699\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__23699\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\
        );

    \I__3111\ : InMux
    port map (
            O => \N__23696\,
            I => \N__23693\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__23693\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23686\
        );

    \I__3108\ : InMux
    port map (
            O => \N__23689\,
            I => \N__23683\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__23686\,
            I => \N__23678\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__23683\,
            I => \N__23678\
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__23678\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__23675\,
            I => \N__23670\
        );

    \I__3103\ : InMux
    port map (
            O => \N__23674\,
            I => \N__23667\
        );

    \I__3102\ : InMux
    port map (
            O => \N__23673\,
            I => \N__23664\
        );

    \I__3101\ : InMux
    port map (
            O => \N__23670\,
            I => \N__23661\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__23667\,
            I => \N__23655\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__23664\,
            I => \N__23655\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__23661\,
            I => \N__23652\
        );

    \I__3097\ : InMux
    port map (
            O => \N__23660\,
            I => \N__23648\
        );

    \I__3096\ : Span4Mux_v
    port map (
            O => \N__23655\,
            I => \N__23645\
        );

    \I__3095\ : Span12Mux_h
    port map (
            O => \N__23652\,
            I => \N__23642\
        );

    \I__3094\ : InMux
    port map (
            O => \N__23651\,
            I => \N__23639\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__23648\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__3092\ : Odrv4
    port map (
            O => \N__23645\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__3091\ : Odrv12
    port map (
            O => \N__23642\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__23639\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__3089\ : InMux
    port map (
            O => \N__23630\,
            I => \N__23627\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__23627\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__23624\,
            I => \N__23620\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23623\,
            I => \N__23617\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23620\,
            I => \N__23614\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__23617\,
            I => \N__23608\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__23614\,
            I => \N__23608\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__23613\,
            I => \N__23605\
        );

    \I__3081\ : Sp12to4
    port map (
            O => \N__23608\,
            I => \N__23602\
        );

    \I__3080\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23599\
        );

    \I__3079\ : Odrv12
    port map (
            O => \N__23602\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__23599\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__3077\ : InMux
    port map (
            O => \N__23594\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__3076\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23588\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__23588\,
            I => \N__23585\
        );

    \I__3074\ : Span12Mux_v
    port map (
            O => \N__23585\,
            I => \N__23582\
        );

    \I__3073\ : Span12Mux_h
    port map (
            O => \N__23582\,
            I => \N__23579\
        );

    \I__3072\ : Odrv12
    port map (
            O => \N__23579\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_12\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__23576\,
            I => \N__23573\
        );

    \I__3070\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23570\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__23570\,
            I => \N__23567\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__23567\,
            I => \current_shift_inst.PI_CTRL.integrator_1_28\
        );

    \I__3067\ : InMux
    port map (
            O => \N__23564\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\
        );

    \I__3066\ : InMux
    port map (
            O => \N__23561\,
            I => \N__23558\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__23558\,
            I => \N__23555\
        );

    \I__3064\ : Span4Mux_v
    port map (
            O => \N__23555\,
            I => \N__23552\
        );

    \I__3063\ : Sp12to4
    port map (
            O => \N__23552\,
            I => \N__23549\
        );

    \I__3062\ : Span12Mux_h
    port map (
            O => \N__23549\,
            I => \N__23546\
        );

    \I__3061\ : Span12Mux_h
    port map (
            O => \N__23546\,
            I => \N__23543\
        );

    \I__3060\ : Odrv12
    port map (
            O => \N__23543\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_13\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__23540\,
            I => \N__23537\
        );

    \I__3058\ : InMux
    port map (
            O => \N__23537\,
            I => \N__23534\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__23534\,
            I => \current_shift_inst.PI_CTRL.integrator_1_29\
        );

    \I__3056\ : InMux
    port map (
            O => \N__23531\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\
        );

    \I__3055\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23525\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__23525\,
            I => \N__23522\
        );

    \I__3053\ : Span4Mux_v
    port map (
            O => \N__23522\,
            I => \N__23519\
        );

    \I__3052\ : Sp12to4
    port map (
            O => \N__23519\,
            I => \N__23516\
        );

    \I__3051\ : Span12Mux_h
    port map (
            O => \N__23516\,
            I => \N__23513\
        );

    \I__3050\ : Span12Mux_h
    port map (
            O => \N__23513\,
            I => \N__23510\
        );

    \I__3049\ : Odrv12
    port map (
            O => \N__23510\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_14\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__23507\,
            I => \N__23504\
        );

    \I__3047\ : InMux
    port map (
            O => \N__23504\,
            I => \N__23501\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__23501\,
            I => \current_shift_inst.PI_CTRL.integrator_1_30\
        );

    \I__3045\ : InMux
    port map (
            O => \N__23498\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\
        );

    \I__3044\ : InMux
    port map (
            O => \N__23495\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__23492\,
            I => \N__23489\
        );

    \I__3042\ : InMux
    port map (
            O => \N__23489\,
            I => \N__23486\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__23486\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\
        );

    \I__3040\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23480\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__23480\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__3038\ : CascadeMux
    port map (
            O => \N__23477\,
            I => \N__23463\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__23476\,
            I => \N__23460\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__23475\,
            I => \N__23457\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__23474\,
            I => \N__23454\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__23473\,
            I => \N__23450\
        );

    \I__3033\ : CascadeMux
    port map (
            O => \N__23472\,
            I => \N__23447\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__23471\,
            I => \N__23444\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__23470\,
            I => \N__23441\
        );

    \I__3030\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23431\
        );

    \I__3029\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23431\
        );

    \I__3028\ : InMux
    port map (
            O => \N__23467\,
            I => \N__23417\
        );

    \I__3027\ : InMux
    port map (
            O => \N__23466\,
            I => \N__23410\
        );

    \I__3026\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23410\
        );

    \I__3025\ : InMux
    port map (
            O => \N__23460\,
            I => \N__23410\
        );

    \I__3024\ : InMux
    port map (
            O => \N__23457\,
            I => \N__23403\
        );

    \I__3023\ : InMux
    port map (
            O => \N__23454\,
            I => \N__23403\
        );

    \I__3022\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23403\
        );

    \I__3021\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23390\
        );

    \I__3020\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23390\
        );

    \I__3019\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23390\
        );

    \I__3018\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23390\
        );

    \I__3017\ : InMux
    port map (
            O => \N__23440\,
            I => \N__23390\
        );

    \I__3016\ : InMux
    port map (
            O => \N__23439\,
            I => \N__23390\
        );

    \I__3015\ : InMux
    port map (
            O => \N__23438\,
            I => \N__23387\
        );

    \I__3014\ : InMux
    port map (
            O => \N__23437\,
            I => \N__23380\
        );

    \I__3013\ : InMux
    port map (
            O => \N__23436\,
            I => \N__23380\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__23431\,
            I => \N__23377\
        );

    \I__3011\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23362\
        );

    \I__3010\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23362\
        );

    \I__3009\ : InMux
    port map (
            O => \N__23428\,
            I => \N__23362\
        );

    \I__3008\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23362\
        );

    \I__3007\ : InMux
    port map (
            O => \N__23426\,
            I => \N__23362\
        );

    \I__3006\ : InMux
    port map (
            O => \N__23425\,
            I => \N__23362\
        );

    \I__3005\ : InMux
    port map (
            O => \N__23424\,
            I => \N__23362\
        );

    \I__3004\ : InMux
    port map (
            O => \N__23423\,
            I => \N__23353\
        );

    \I__3003\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23353\
        );

    \I__3002\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23353\
        );

    \I__3001\ : InMux
    port map (
            O => \N__23420\,
            I => \N__23353\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__23417\,
            I => \N__23350\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__23410\,
            I => \N__23345\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__23403\,
            I => \N__23345\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__23390\,
            I => \N__23340\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__23387\,
            I => \N__23340\
        );

    \I__2995\ : InMux
    port map (
            O => \N__23386\,
            I => \N__23335\
        );

    \I__2994\ : InMux
    port map (
            O => \N__23385\,
            I => \N__23335\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__23380\,
            I => \N__23330\
        );

    \I__2992\ : Span4Mux_h
    port map (
            O => \N__23377\,
            I => \N__23330\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__23362\,
            I => \N__23321\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__23353\,
            I => \N__23321\
        );

    \I__2989\ : Span4Mux_h
    port map (
            O => \N__23350\,
            I => \N__23321\
        );

    \I__2988\ : Span4Mux_v
    port map (
            O => \N__23345\,
            I => \N__23321\
        );

    \I__2987\ : Span4Mux_v
    port map (
            O => \N__23340\,
            I => \N__23318\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__23335\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2985\ : Odrv4
    port map (
            O => \N__23330\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__23321\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2983\ : Odrv4
    port map (
            O => \N__23318\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2982\ : InMux
    port map (
            O => \N__23309\,
            I => \N__23306\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__23306\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__2980\ : InMux
    port map (
            O => \N__23303\,
            I => \N__23300\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__23300\,
            I => \N__23297\
        );

    \I__2978\ : Span4Mux_h
    port map (
            O => \N__23297\,
            I => \N__23294\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__23294\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\
        );

    \I__2976\ : InMux
    port map (
            O => \N__23291\,
            I => \N__23288\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__23288\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__23285\,
            I => \N__23265\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__23284\,
            I => \N__23259\
        );

    \I__2972\ : InMux
    port map (
            O => \N__23283\,
            I => \N__23245\
        );

    \I__2971\ : InMux
    port map (
            O => \N__23282\,
            I => \N__23245\
        );

    \I__2970\ : InMux
    port map (
            O => \N__23281\,
            I => \N__23245\
        );

    \I__2969\ : InMux
    port map (
            O => \N__23280\,
            I => \N__23245\
        );

    \I__2968\ : InMux
    port map (
            O => \N__23279\,
            I => \N__23245\
        );

    \I__2967\ : InMux
    port map (
            O => \N__23278\,
            I => \N__23245\
        );

    \I__2966\ : InMux
    port map (
            O => \N__23277\,
            I => \N__23240\
        );

    \I__2965\ : InMux
    port map (
            O => \N__23276\,
            I => \N__23240\
        );

    \I__2964\ : InMux
    port map (
            O => \N__23275\,
            I => \N__23233\
        );

    \I__2963\ : InMux
    port map (
            O => \N__23274\,
            I => \N__23233\
        );

    \I__2962\ : InMux
    port map (
            O => \N__23273\,
            I => \N__23233\
        );

    \I__2961\ : InMux
    port map (
            O => \N__23272\,
            I => \N__23226\
        );

    \I__2960\ : InMux
    port map (
            O => \N__23271\,
            I => \N__23226\
        );

    \I__2959\ : InMux
    port map (
            O => \N__23270\,
            I => \N__23226\
        );

    \I__2958\ : InMux
    port map (
            O => \N__23269\,
            I => \N__23217\
        );

    \I__2957\ : InMux
    port map (
            O => \N__23268\,
            I => \N__23214\
        );

    \I__2956\ : InMux
    port map (
            O => \N__23265\,
            I => \N__23209\
        );

    \I__2955\ : InMux
    port map (
            O => \N__23264\,
            I => \N__23209\
        );

    \I__2954\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23200\
        );

    \I__2953\ : InMux
    port map (
            O => \N__23262\,
            I => \N__23200\
        );

    \I__2952\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23200\
        );

    \I__2951\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23200\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__23245\,
            I => \N__23197\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__23240\,
            I => \N__23192\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__23233\,
            I => \N__23192\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__23226\,
            I => \N__23189\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__23225\,
            I => \N__23186\
        );

    \I__2945\ : CascadeMux
    port map (
            O => \N__23224\,
            I => \N__23183\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__23223\,
            I => \N__23178\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__23222\,
            I => \N__23175\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__23221\,
            I => \N__23172\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__23220\,
            I => \N__23169\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__23217\,
            I => \N__23165\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__23214\,
            I => \N__23162\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__23209\,
            I => \N__23159\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__23200\,
            I => \N__23150\
        );

    \I__2936\ : Span4Mux_h
    port map (
            O => \N__23197\,
            I => \N__23150\
        );

    \I__2935\ : Span4Mux_h
    port map (
            O => \N__23192\,
            I => \N__23150\
        );

    \I__2934\ : Span4Mux_v
    port map (
            O => \N__23189\,
            I => \N__23150\
        );

    \I__2933\ : InMux
    port map (
            O => \N__23186\,
            I => \N__23145\
        );

    \I__2932\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23145\
        );

    \I__2931\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23130\
        );

    \I__2930\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23130\
        );

    \I__2929\ : InMux
    port map (
            O => \N__23178\,
            I => \N__23130\
        );

    \I__2928\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23130\
        );

    \I__2927\ : InMux
    port map (
            O => \N__23172\,
            I => \N__23130\
        );

    \I__2926\ : InMux
    port map (
            O => \N__23169\,
            I => \N__23130\
        );

    \I__2925\ : InMux
    port map (
            O => \N__23168\,
            I => \N__23130\
        );

    \I__2924\ : Span4Mux_h
    port map (
            O => \N__23165\,
            I => \N__23127\
        );

    \I__2923\ : Span4Mux_v
    port map (
            O => \N__23162\,
            I => \N__23124\
        );

    \I__2922\ : Span4Mux_v
    port map (
            O => \N__23159\,
            I => \N__23119\
        );

    \I__2921\ : Span4Mux_v
    port map (
            O => \N__23150\,
            I => \N__23119\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__23145\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__23130\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2918\ : Odrv4
    port map (
            O => \N__23127\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__23124\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2916\ : Odrv4
    port map (
            O => \N__23119\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2915\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23105\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__23105\,
            I => \N__23102\
        );

    \I__2913\ : Span12Mux_v
    port map (
            O => \N__23102\,
            I => \N__23099\
        );

    \I__2912\ : Span12Mux_h
    port map (
            O => \N__23099\,
            I => \N__23096\
        );

    \I__2911\ : Odrv12
    port map (
            O => \N__23096\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_4\
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__23093\,
            I => \N__23090\
        );

    \I__2909\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23087\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__23087\,
            I => \N__23084\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__23084\,
            I => \current_shift_inst.PI_CTRL.integrator_1_20\
        );

    \I__2906\ : InMux
    port map (
            O => \N__23081\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\
        );

    \I__2905\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23075\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__23075\,
            I => \N__23072\
        );

    \I__2903\ : Span4Mux_h
    port map (
            O => \N__23072\,
            I => \N__23069\
        );

    \I__2902\ : Sp12to4
    port map (
            O => \N__23069\,
            I => \N__23066\
        );

    \I__2901\ : Span12Mux_v
    port map (
            O => \N__23066\,
            I => \N__23063\
        );

    \I__2900\ : Span12Mux_h
    port map (
            O => \N__23063\,
            I => \N__23060\
        );

    \I__2899\ : Odrv12
    port map (
            O => \N__23060\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_5\
        );

    \I__2898\ : CascadeMux
    port map (
            O => \N__23057\,
            I => \N__23054\
        );

    \I__2897\ : InMux
    port map (
            O => \N__23054\,
            I => \N__23051\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__23051\,
            I => \N__23048\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__23048\,
            I => \current_shift_inst.PI_CTRL.integrator_1_21\
        );

    \I__2894\ : InMux
    port map (
            O => \N__23045\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\
        );

    \I__2893\ : InMux
    port map (
            O => \N__23042\,
            I => \N__23039\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__23039\,
            I => \N__23036\
        );

    \I__2891\ : Span4Mux_v
    port map (
            O => \N__23036\,
            I => \N__23033\
        );

    \I__2890\ : Sp12to4
    port map (
            O => \N__23033\,
            I => \N__23030\
        );

    \I__2889\ : Span12Mux_h
    port map (
            O => \N__23030\,
            I => \N__23027\
        );

    \I__2888\ : Span12Mux_h
    port map (
            O => \N__23027\,
            I => \N__23024\
        );

    \I__2887\ : Odrv12
    port map (
            O => \N__23024\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_6\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__23021\,
            I => \N__23018\
        );

    \I__2885\ : InMux
    port map (
            O => \N__23018\,
            I => \N__23015\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__23015\,
            I => \current_shift_inst.PI_CTRL.integrator_1_22\
        );

    \I__2883\ : InMux
    port map (
            O => \N__23012\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\
        );

    \I__2882\ : InMux
    port map (
            O => \N__23009\,
            I => \N__23006\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__23006\,
            I => \N__23003\
        );

    \I__2880\ : Span4Mux_v
    port map (
            O => \N__23003\,
            I => \N__23000\
        );

    \I__2879\ : Sp12to4
    port map (
            O => \N__23000\,
            I => \N__22997\
        );

    \I__2878\ : Span12Mux_h
    port map (
            O => \N__22997\,
            I => \N__22994\
        );

    \I__2877\ : Span12Mux_v
    port map (
            O => \N__22994\,
            I => \N__22991\
        );

    \I__2876\ : Odrv12
    port map (
            O => \N__22991\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_7\
        );

    \I__2875\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22985\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__22985\,
            I => \current_shift_inst.PI_CTRL.integrator_1_23\
        );

    \I__2873\ : InMux
    port map (
            O => \N__22982\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__22979\,
            I => \N__22976\
        );

    \I__2871\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22973\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__22973\,
            I => \N__22970\
        );

    \I__2869\ : Span4Mux_v
    port map (
            O => \N__22970\,
            I => \N__22967\
        );

    \I__2868\ : Sp12to4
    port map (
            O => \N__22967\,
            I => \N__22964\
        );

    \I__2867\ : Span12Mux_h
    port map (
            O => \N__22964\,
            I => \N__22961\
        );

    \I__2866\ : Span12Mux_h
    port map (
            O => \N__22961\,
            I => \N__22958\
        );

    \I__2865\ : Odrv12
    port map (
            O => \N__22958\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_8\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__22955\,
            I => \N__22952\
        );

    \I__2863\ : InMux
    port map (
            O => \N__22952\,
            I => \N__22949\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__22949\,
            I => \current_shift_inst.PI_CTRL.integrator_1_24\
        );

    \I__2861\ : InMux
    port map (
            O => \N__22946\,
            I => \bfn_5_15_0_\
        );

    \I__2860\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22940\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__22940\,
            I => \N__22937\
        );

    \I__2858\ : Span4Mux_h
    port map (
            O => \N__22937\,
            I => \N__22934\
        );

    \I__2857\ : Sp12to4
    port map (
            O => \N__22934\,
            I => \N__22931\
        );

    \I__2856\ : Span12Mux_v
    port map (
            O => \N__22931\,
            I => \N__22928\
        );

    \I__2855\ : Span12Mux_h
    port map (
            O => \N__22928\,
            I => \N__22925\
        );

    \I__2854\ : Odrv12
    port map (
            O => \N__22925\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_9\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__22922\,
            I => \N__22919\
        );

    \I__2852\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22916\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__22916\,
            I => \current_shift_inst.PI_CTRL.integrator_1_25\
        );

    \I__2850\ : InMux
    port map (
            O => \N__22913\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__22910\,
            I => \N__22907\
        );

    \I__2848\ : InMux
    port map (
            O => \N__22907\,
            I => \N__22904\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__22904\,
            I => \N__22901\
        );

    \I__2846\ : Span4Mux_v
    port map (
            O => \N__22901\,
            I => \N__22898\
        );

    \I__2845\ : Sp12to4
    port map (
            O => \N__22898\,
            I => \N__22895\
        );

    \I__2844\ : Span12Mux_h
    port map (
            O => \N__22895\,
            I => \N__22892\
        );

    \I__2843\ : Span12Mux_h
    port map (
            O => \N__22892\,
            I => \N__22889\
        );

    \I__2842\ : Odrv12
    port map (
            O => \N__22889\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_10\
        );

    \I__2841\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22883\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__22883\,
            I => \current_shift_inst.PI_CTRL.integrator_1_26\
        );

    \I__2839\ : InMux
    port map (
            O => \N__22880\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\
        );

    \I__2838\ : InMux
    port map (
            O => \N__22877\,
            I => \N__22874\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__22874\,
            I => \N__22871\
        );

    \I__2836\ : Span12Mux_h
    port map (
            O => \N__22871\,
            I => \N__22868\
        );

    \I__2835\ : Span12Mux_h
    port map (
            O => \N__22868\,
            I => \N__22865\
        );

    \I__2834\ : Odrv12
    port map (
            O => \N__22865\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_11\
        );

    \I__2833\ : CascadeMux
    port map (
            O => \N__22862\,
            I => \N__22859\
        );

    \I__2832\ : InMux
    port map (
            O => \N__22859\,
            I => \N__22856\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__22856\,
            I => \current_shift_inst.PI_CTRL.integrator_1_27\
        );

    \I__2830\ : InMux
    port map (
            O => \N__22853\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\
        );

    \I__2829\ : InMux
    port map (
            O => \N__22850\,
            I => \N__22847\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__22847\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__2827\ : InMux
    port map (
            O => \N__22844\,
            I => \N__22841\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__22841\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__2825\ : CascadeMux
    port map (
            O => \N__22838\,
            I => \N__22835\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22832\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__22832\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__2822\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22826\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__22826\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__2820\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22820\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__22820\,
            I => \N__22817\
        );

    \I__2818\ : Span4Mux_h
    port map (
            O => \N__22817\,
            I => \N__22814\
        );

    \I__2817\ : Span4Mux_h
    port map (
            O => \N__22814\,
            I => \N__22811\
        );

    \I__2816\ : Odrv4
    port map (
            O => \N__22811\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_15\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__22808\,
            I => \N__22805\
        );

    \I__2814\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22802\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__22802\,
            I => \N__22799\
        );

    \I__2812\ : Span4Mux_v
    port map (
            O => \N__22799\,
            I => \N__22796\
        );

    \I__2811\ : Sp12to4
    port map (
            O => \N__22796\,
            I => \N__22793\
        );

    \I__2810\ : Span12Mux_h
    port map (
            O => \N__22793\,
            I => \N__22790\
        );

    \I__2809\ : Span12Mux_h
    port map (
            O => \N__22790\,
            I => \N__22787\
        );

    \I__2808\ : Odrv12
    port map (
            O => \N__22787\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_0\
        );

    \I__2807\ : CascadeMux
    port map (
            O => \N__22784\,
            I => \N__22781\
        );

    \I__2806\ : InMux
    port map (
            O => \N__22781\,
            I => \N__22778\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__22778\,
            I => \N__22775\
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__22775\,
            I => \current_shift_inst.PI_CTRL.integrator_1_16\
        );

    \I__2803\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22769\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__22769\,
            I => \N__22766\
        );

    \I__2801\ : Span4Mux_h
    port map (
            O => \N__22766\,
            I => \N__22763\
        );

    \I__2800\ : Sp12to4
    port map (
            O => \N__22763\,
            I => \N__22760\
        );

    \I__2799\ : Span12Mux_v
    port map (
            O => \N__22760\,
            I => \N__22757\
        );

    \I__2798\ : Span12Mux_h
    port map (
            O => \N__22757\,
            I => \N__22754\
        );

    \I__2797\ : Odrv12
    port map (
            O => \N__22754\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_1\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__22751\,
            I => \N__22748\
        );

    \I__2795\ : InMux
    port map (
            O => \N__22748\,
            I => \N__22745\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__22745\,
            I => \N__22742\
        );

    \I__2793\ : Span4Mux_h
    port map (
            O => \N__22742\,
            I => \N__22739\
        );

    \I__2792\ : Span4Mux_h
    port map (
            O => \N__22739\,
            I => \N__22736\
        );

    \I__2791\ : Odrv4
    port map (
            O => \N__22736\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_16\
        );

    \I__2790\ : CascadeMux
    port map (
            O => \N__22733\,
            I => \N__22730\
        );

    \I__2789\ : InMux
    port map (
            O => \N__22730\,
            I => \N__22727\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__22727\,
            I => \current_shift_inst.PI_CTRL.integrator_1_17\
        );

    \I__2787\ : InMux
    port map (
            O => \N__22724\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\
        );

    \I__2786\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22718\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__22718\,
            I => \N__22715\
        );

    \I__2784\ : Span4Mux_v
    port map (
            O => \N__22715\,
            I => \N__22712\
        );

    \I__2783\ : Sp12to4
    port map (
            O => \N__22712\,
            I => \N__22709\
        );

    \I__2782\ : Span12Mux_h
    port map (
            O => \N__22709\,
            I => \N__22706\
        );

    \I__2781\ : Span12Mux_v
    port map (
            O => \N__22706\,
            I => \N__22703\
        );

    \I__2780\ : Odrv12
    port map (
            O => \N__22703\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_2\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__22700\,
            I => \N__22697\
        );

    \I__2778\ : InMux
    port map (
            O => \N__22697\,
            I => \N__22694\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__22694\,
            I => \N__22691\
        );

    \I__2776\ : Span4Mux_h
    port map (
            O => \N__22691\,
            I => \N__22688\
        );

    \I__2775\ : Span4Mux_h
    port map (
            O => \N__22688\,
            I => \N__22685\
        );

    \I__2774\ : Odrv4
    port map (
            O => \N__22685\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_17\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__22682\,
            I => \N__22679\
        );

    \I__2772\ : InMux
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__22676\,
            I => \current_shift_inst.PI_CTRL.integrator_1_18\
        );

    \I__2770\ : InMux
    port map (
            O => \N__22673\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\
        );

    \I__2769\ : InMux
    port map (
            O => \N__22670\,
            I => \N__22667\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__22667\,
            I => \N__22664\
        );

    \I__2767\ : Span12Mux_h
    port map (
            O => \N__22664\,
            I => \N__22661\
        );

    \I__2766\ : Span12Mux_v
    port map (
            O => \N__22661\,
            I => \N__22658\
        );

    \I__2765\ : Span12Mux_h
    port map (
            O => \N__22658\,
            I => \N__22655\
        );

    \I__2764\ : Odrv12
    port map (
            O => \N__22655\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_3\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__22652\,
            I => \N__22649\
        );

    \I__2762\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22646\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__22646\,
            I => \N__22643\
        );

    \I__2760\ : Span12Mux_h
    port map (
            O => \N__22643\,
            I => \N__22640\
        );

    \I__2759\ : Odrv12
    port map (
            O => \N__22640\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_18\
        );

    \I__2758\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22634\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__22634\,
            I => \current_shift_inst.PI_CTRL.integrator_1_19\
        );

    \I__2756\ : InMux
    port map (
            O => \N__22631\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\
        );

    \I__2755\ : CascadeMux
    port map (
            O => \N__22628\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\
        );

    \I__2754\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22622\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__22622\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2752\ : InMux
    port map (
            O => \N__22619\,
            I => \N__22616\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__22616\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__2750\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22610\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__22610\,
            I => \N__22607\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__22607\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__2747\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22601\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__22601\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__22598\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_\
        );

    \I__2744\ : InMux
    port map (
            O => \N__22595\,
            I => \N__22592\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__22592\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2742\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22585\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22588\,
            I => \N__22582\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__22585\,
            I => \N__22579\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__22582\,
            I => \N__22576\
        );

    \I__2738\ : Span4Mux_h
    port map (
            O => \N__22579\,
            I => \N__22573\
        );

    \I__2737\ : Odrv4
    port map (
            O => \N__22576\,
            I => pwm_duty_input_0
        );

    \I__2736\ : Odrv4
    port map (
            O => \N__22573\,
            I => pwm_duty_input_0
        );

    \I__2735\ : InMux
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__22565\,
            I => \N__22562\
        );

    \I__2733\ : Odrv12
    port map (
            O => \N__22562\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2732\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22555\
        );

    \I__2731\ : InMux
    port map (
            O => \N__22558\,
            I => \N__22552\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__22555\,
            I => \N__22549\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__22552\,
            I => \N__22546\
        );

    \I__2728\ : Span4Mux_h
    port map (
            O => \N__22549\,
            I => \N__22543\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__22546\,
            I => pwm_duty_input_1
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__22543\,
            I => pwm_duty_input_1
        );

    \I__2725\ : InMux
    port map (
            O => \N__22538\,
            I => \N__22535\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__22535\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__2723\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22529\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__22529\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__2721\ : CascadeMux
    port map (
            O => \N__22526\,
            I => \N__22523\
        );

    \I__2720\ : InMux
    port map (
            O => \N__22523\,
            I => \N__22520\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__22520\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__2718\ : CascadeMux
    port map (
            O => \N__22517\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\
        );

    \I__2717\ : InMux
    port map (
            O => \N__22514\,
            I => \N__22511\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__22511\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__2715\ : InMux
    port map (
            O => \N__22508\,
            I => \N__22505\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__22505\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__22502\,
            I => \N__22499\
        );

    \I__2712\ : InMux
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__22496\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2710\ : InMux
    port map (
            O => \N__22493\,
            I => \N__22490\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__22490\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__2708\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22484\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__22484\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__22481\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\
        );

    \I__2705\ : InMux
    port map (
            O => \N__22478\,
            I => \N__22475\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__22475\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\
        );

    \I__2703\ : InMux
    port map (
            O => \N__22472\,
            I => \N__22469\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__22469\,
            I => \current_shift_inst.PI_CTRL.N_77\
        );

    \I__2701\ : InMux
    port map (
            O => \N__22466\,
            I => \N__22463\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__22463\,
            I => \N__22460\
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__22460\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__22457\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__22454\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\
        );

    \I__2696\ : InMux
    port map (
            O => \N__22451\,
            I => \N__22448\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__22448\,
            I => \N__22445\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__22445\,
            I => \current_shift_inst.PI_CTRL.N_44\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__22442\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__2692\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22436\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__22436\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__22433\,
            I => \N__22430\
        );

    \I__2689\ : InMux
    port map (
            O => \N__22430\,
            I => \N__22427\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__22427\,
            I => \N__22424\
        );

    \I__2687\ : Odrv12
    port map (
            O => \N__22424\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__2686\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22418\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__22418\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__22415\,
            I => \N__22412\
        );

    \I__2683\ : InMux
    port map (
            O => \N__22412\,
            I => \N__22409\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__22409\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__2681\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__22403\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__2679\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22397\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__22397\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__22394\,
            I => \N__22391\
        );

    \I__2676\ : InMux
    port map (
            O => \N__22391\,
            I => \N__22388\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__22388\,
            I => \N__22385\
        );

    \I__2674\ : Span4Mux_h
    port map (
            O => \N__22385\,
            I => \N__22382\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__22382\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__2672\ : InMux
    port map (
            O => \N__22379\,
            I => \N__22376\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__22376\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__22373\,
            I => \N__22370\
        );

    \I__2669\ : InMux
    port map (
            O => \N__22370\,
            I => \N__22367\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__2667\ : Span4Mux_h
    port map (
            O => \N__22364\,
            I => \N__22361\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__22361\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\
        );

    \I__2665\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__22355\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__2663\ : InMux
    port map (
            O => \N__22352\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\
        );

    \I__2662\ : InMux
    port map (
            O => \N__22349\,
            I => \bfn_4_15_0_\
        );

    \I__2661\ : InMux
    port map (
            O => \N__22346\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__2660\ : InMux
    port map (
            O => \N__22343\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__2659\ : InMux
    port map (
            O => \N__22340\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__2658\ : InMux
    port map (
            O => \N__22337\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__2657\ : InMux
    port map (
            O => \N__22334\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__2656\ : InMux
    port map (
            O => \N__22331\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__2654\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__22319\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__2650\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__2648\ : Odrv4
    port map (
            O => \N__22307\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__2647\ : InMux
    port map (
            O => \N__22304\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\
        );

    \I__2646\ : InMux
    port map (
            O => \N__22301\,
            I => \bfn_4_14_0_\
        );

    \I__2645\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__22295\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__2643\ : InMux
    port map (
            O => \N__22292\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__22289\,
            I => \N__22286\
        );

    \I__2641\ : InMux
    port map (
            O => \N__22286\,
            I => \N__22283\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__22283\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__2639\ : InMux
    port map (
            O => \N__22280\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__2638\ : InMux
    port map (
            O => \N__22277\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__2637\ : InMux
    port map (
            O => \N__22274\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__2636\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22268\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__22268\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__2634\ : InMux
    port map (
            O => \N__22265\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__22262\,
            I => \N__22259\
        );

    \I__2632\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22256\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__22256\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__2630\ : InMux
    port map (
            O => \N__22253\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__22250\,
            I => \N__22247\
        );

    \I__2628\ : InMux
    port map (
            O => \N__22247\,
            I => \N__22244\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__22244\,
            I => \N__22241\
        );

    \I__2626\ : Span4Mux_h
    port map (
            O => \N__22241\,
            I => \N__22238\
        );

    \I__2625\ : Span4Mux_h
    port map (
            O => \N__22238\,
            I => \N__22235\
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__22235\,
            I => \current_shift_inst.PI_CTRL.integrator_1_8\
        );

    \I__2623\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22229\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__22229\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__2621\ : InMux
    port map (
            O => \N__22226\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__22223\,
            I => \N__22220\
        );

    \I__2619\ : InMux
    port map (
            O => \N__22220\,
            I => \N__22217\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__22217\,
            I => \N__22214\
        );

    \I__2617\ : Span4Mux_v
    port map (
            O => \N__22214\,
            I => \N__22211\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__22211\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__22208\,
            I => \N__22205\
        );

    \I__2614\ : InMux
    port map (
            O => \N__22205\,
            I => \N__22202\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__22202\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__2612\ : InMux
    port map (
            O => \N__22199\,
            I => \bfn_4_13_0_\
        );

    \I__2611\ : CascadeMux
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__2610\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__22184\,
            I => \current_shift_inst.PI_CTRL.integrator_1_10\
        );

    \I__2606\ : InMux
    port map (
            O => \N__22181\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__22178\,
            I => \N__22175\
        );

    \I__2604\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__22172\,
            I => \N__22169\
        );

    \I__2602\ : Span4Mux_v
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__2601\ : Span4Mux_h
    port map (
            O => \N__22166\,
            I => \N__22163\
        );

    \I__2600\ : Odrv4
    port map (
            O => \N__22163\,
            I => \current_shift_inst.PI_CTRL.integrator_1_11\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__22160\,
            I => \N__22157\
        );

    \I__2598\ : InMux
    port map (
            O => \N__22157\,
            I => \N__22154\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__22154\,
            I => \N__22151\
        );

    \I__2596\ : Span4Mux_h
    port map (
            O => \N__22151\,
            I => \N__22148\
        );

    \I__2595\ : Odrv4
    port map (
            O => \N__22148\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__2594\ : InMux
    port map (
            O => \N__22145\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__2593\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__22139\,
            I => \N__22136\
        );

    \I__2591\ : Span4Mux_v
    port map (
            O => \N__22136\,
            I => \N__22133\
        );

    \I__2590\ : Odrv4
    port map (
            O => \N__22133\,
            I => \current_shift_inst.PI_CTRL.integrator_1_12\
        );

    \I__2589\ : InMux
    port map (
            O => \N__22130\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__22127\,
            I => \N__22124\
        );

    \I__2587\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22121\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__22121\,
            I => \N__22118\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__22118\,
            I => \N__22115\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__22115\,
            I => \current_shift_inst.PI_CTRL.integrator_1_13\
        );

    \I__2583\ : InMux
    port map (
            O => \N__22112\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__22109\,
            I => \N__22106\
        );

    \I__2581\ : InMux
    port map (
            O => \N__22106\,
            I => \N__22103\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__22103\,
            I => \N__22100\
        );

    \I__2579\ : Span4Mux_h
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__2578\ : Odrv4
    port map (
            O => \N__22097\,
            I => \current_shift_inst.PI_CTRL.integrator_1_14\
        );

    \I__2577\ : InMux
    port map (
            O => \N__22094\,
            I => \N__22091\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__22091\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__2575\ : InMux
    port map (
            O => \N__22088\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__2574\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22082\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__22082\,
            I => \N__22079\
        );

    \I__2572\ : Span4Mux_h
    port map (
            O => \N__22079\,
            I => \N__22076\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__22076\,
            I => \current_shift_inst.PI_CTRL.integrator_1_15\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__22073\,
            I => \N__22070\
        );

    \I__2569\ : InMux
    port map (
            O => \N__22070\,
            I => \N__22067\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__22067\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__2567\ : InMux
    port map (
            O => \N__22064\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__2566\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22058\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__22058\,
            I => \N__22053\
        );

    \I__2564\ : InMux
    port map (
            O => \N__22057\,
            I => \N__22048\
        );

    \I__2563\ : InMux
    port map (
            O => \N__22056\,
            I => \N__22048\
        );

    \I__2562\ : Span4Mux_s3_h
    port map (
            O => \N__22053\,
            I => \N__22045\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__22048\,
            I => pwm_duty_input_7
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__22045\,
            I => pwm_duty_input_7
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__22040\,
            I => \N__22036\
        );

    \I__2558\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22033\
        );

    \I__2557\ : InMux
    port map (
            O => \N__22036\,
            I => \N__22030\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__22033\,
            I => \N__22025\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__22030\,
            I => \N__22025\
        );

    \I__2554\ : Span4Mux_v
    port map (
            O => \N__22025\,
            I => \N__22022\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__22022\,
            I => \current_shift_inst.PI_CTRL.un1_integrator\
        );

    \I__2552\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22016\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__22016\,
            I => \N__22013\
        );

    \I__2550\ : Span4Mux_v
    port map (
            O => \N__22013\,
            I => \N__22010\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__22010\,
            I => \current_shift_inst.PI_CTRL.integrator_1_2\
        );

    \I__2548\ : InMux
    port map (
            O => \N__22007\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__2547\ : CascadeMux
    port map (
            O => \N__22004\,
            I => \N__22001\
        );

    \I__2546\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__21995\,
            I => \N__21992\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__21992\,
            I => \current_shift_inst.PI_CTRL.integrator_1_3\
        );

    \I__2542\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21986\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__21986\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__2540\ : InMux
    port map (
            O => \N__21983\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__2539\ : InMux
    port map (
            O => \N__21980\,
            I => \N__21977\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__21977\,
            I => \N__21974\
        );

    \I__2537\ : Span4Mux_v
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__21971\,
            I => \current_shift_inst.PI_CTRL.integrator_1_4\
        );

    \I__2535\ : InMux
    port map (
            O => \N__21968\,
            I => \N__21965\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__21965\,
            I => \N__21962\
        );

    \I__2533\ : Span4Mux_h
    port map (
            O => \N__21962\,
            I => \N__21959\
        );

    \I__2532\ : Odrv4
    port map (
            O => \N__21959\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__2531\ : InMux
    port map (
            O => \N__21956\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__2530\ : CascadeMux
    port map (
            O => \N__21953\,
            I => \N__21950\
        );

    \I__2529\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__2527\ : Span4Mux_v
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__21941\,
            I => \current_shift_inst.PI_CTRL.integrator_1_5\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__2524\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21932\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__2522\ : Span4Mux_v
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__2521\ : Odrv4
    port map (
            O => \N__21926\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__2520\ : InMux
    port map (
            O => \N__21923\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__21920\,
            I => \N__21917\
        );

    \I__2518\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21914\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__21914\,
            I => \N__21911\
        );

    \I__2516\ : Span4Mux_v
    port map (
            O => \N__21911\,
            I => \N__21908\
        );

    \I__2515\ : Odrv4
    port map (
            O => \N__21908\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__2514\ : InMux
    port map (
            O => \N__21905\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__21902\,
            I => \N__21899\
        );

    \I__2512\ : InMux
    port map (
            O => \N__21899\,
            I => \N__21896\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__21896\,
            I => \N__21893\
        );

    \I__2510\ : Span4Mux_h
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__21890\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__2508\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21884\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__21884\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__2506\ : InMux
    port map (
            O => \N__21881\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__21878\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\
        );

    \I__2504\ : InMux
    port map (
            O => \N__21875\,
            I => \N__21872\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__21872\,
            I => \N__21869\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__21869\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\
        );

    \I__2501\ : InMux
    port map (
            O => \N__21866\,
            I => \N__21863\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__21863\,
            I => \N__21860\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__21860\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__21857\,
            I => \current_shift_inst.PI_CTRL.N_98_cascade_\
        );

    \I__2497\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21851\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__21851\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__2495\ : CascadeMux
    port map (
            O => \N__21848\,
            I => \current_shift_inst.PI_CTRL.N_96_cascade_\
        );

    \I__2494\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21841\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__21844\,
            I => \N__21838\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__21841\,
            I => \N__21834\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21838\,
            I => \N__21829\
        );

    \I__2490\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21829\
        );

    \I__2489\ : Span4Mux_s3_h
    port map (
            O => \N__21834\,
            I => \N__21826\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__21829\,
            I => pwm_duty_input_6
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__21826\,
            I => pwm_duty_input_6
        );

    \I__2486\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21818\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__21818\,
            I => \N__21815\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__21815\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__21812\,
            I => \N__21809\
        );

    \I__2482\ : InMux
    port map (
            O => \N__21809\,
            I => \N__21805\
        );

    \I__2481\ : InMux
    port map (
            O => \N__21808\,
            I => \N__21802\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__21805\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__21802\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__2477\ : InMux
    port map (
            O => \N__21794\,
            I => \N__21789\
        );

    \I__2476\ : InMux
    port map (
            O => \N__21793\,
            I => \N__21786\
        );

    \I__2475\ : InMux
    port map (
            O => \N__21792\,
            I => \N__21783\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__21789\,
            I => \N__21780\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__21786\,
            I => \N__21777\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__21783\,
            I => \N__21774\
        );

    \I__2471\ : Span4Mux_v
    port map (
            O => \N__21780\,
            I => \N__21767\
        );

    \I__2470\ : Span4Mux_v
    port map (
            O => \N__21777\,
            I => \N__21767\
        );

    \I__2469\ : Span4Mux_s3_h
    port map (
            O => \N__21774\,
            I => \N__21767\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__21767\,
            I => pwm_duty_input_4
        );

    \I__2467\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21760\
        );

    \I__2466\ : InMux
    port map (
            O => \N__21763\,
            I => \N__21757\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__21760\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__21757\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__2463\ : InMux
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__21749\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__2461\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21741\
        );

    \I__2460\ : InMux
    port map (
            O => \N__21745\,
            I => \N__21738\
        );

    \I__2459\ : InMux
    port map (
            O => \N__21744\,
            I => \N__21735\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__21741\,
            I => \N__21732\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__21738\,
            I => \N__21727\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__21735\,
            I => \N__21727\
        );

    \I__2455\ : Span4Mux_s3_h
    port map (
            O => \N__21732\,
            I => \N__21724\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__21727\,
            I => pwm_duty_input_3
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__21724\,
            I => pwm_duty_input_3
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__21719\,
            I => \N__21715\
        );

    \I__2451\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21712\
        );

    \I__2450\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21709\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__21712\,
            I => \N__21705\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__21709\,
            I => \N__21702\
        );

    \I__2447\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21699\
        );

    \I__2446\ : Span4Mux_s3_h
    port map (
            O => \N__21705\,
            I => \N__21696\
        );

    \I__2445\ : Odrv12
    port map (
            O => \N__21702\,
            I => pwm_duty_input_5
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__21699\,
            I => pwm_duty_input_5
        );

    \I__2443\ : Odrv4
    port map (
            O => \N__21696\,
            I => pwm_duty_input_5
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__21689\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11_cascade_\
        );

    \I__2441\ : CascadeMux
    port map (
            O => \N__21686\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__21683\,
            I => \current_shift_inst.PI_CTRL.N_31_cascade_\
        );

    \I__2439\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__21677\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4\
        );

    \I__2437\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21670\
        );

    \I__2436\ : InMux
    port map (
            O => \N__21673\,
            I => \N__21667\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__21670\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__21667\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__21662\,
            I => \N__21659\
        );

    \I__2432\ : InMux
    port map (
            O => \N__21659\,
            I => \N__21656\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__21656\,
            I => \pwm_generator_inst.threshold_9\
        );

    \I__2430\ : InMux
    port map (
            O => \N__21653\,
            I => \N__21650\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__21650\,
            I => \N__21646\
        );

    \I__2428\ : InMux
    port map (
            O => \N__21649\,
            I => \N__21642\
        );

    \I__2427\ : Span4Mux_h
    port map (
            O => \N__21646\,
            I => \N__21639\
        );

    \I__2426\ : InMux
    port map (
            O => \N__21645\,
            I => \N__21636\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__21642\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2424\ : Odrv4
    port map (
            O => \N__21639\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__21636\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2422\ : InMux
    port map (
            O => \N__21629\,
            I => \N__21626\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__21626\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2420\ : InMux
    port map (
            O => \N__21623\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2419\ : IoInMux
    port map (
            O => \N__21620\,
            I => \N__21617\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__21617\,
            I => \N__21614\
        );

    \I__2417\ : Span4Mux_s2_v
    port map (
            O => \N__21614\,
            I => \N__21611\
        );

    \I__2416\ : Sp12to4
    port map (
            O => \N__21611\,
            I => \N__21608\
        );

    \I__2415\ : Span12Mux_s10_h
    port map (
            O => \N__21608\,
            I => \N__21605\
        );

    \I__2414\ : Span12Mux_h
    port map (
            O => \N__21605\,
            I => \N__21602\
        );

    \I__2413\ : Span12Mux_v
    port map (
            O => \N__21602\,
            I => \N__21599\
        );

    \I__2412\ : Odrv12
    port map (
            O => \N__21599\,
            I => pwm_output_c
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__21596\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__2410\ : InMux
    port map (
            O => \N__21593\,
            I => \N__21573\
        );

    \I__2409\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21573\
        );

    \I__2408\ : InMux
    port map (
            O => \N__21591\,
            I => \N__21573\
        );

    \I__2407\ : InMux
    port map (
            O => \N__21590\,
            I => \N__21573\
        );

    \I__2406\ : InMux
    port map (
            O => \N__21589\,
            I => \N__21573\
        );

    \I__2405\ : InMux
    port map (
            O => \N__21588\,
            I => \N__21564\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21587\,
            I => \N__21564\
        );

    \I__2403\ : InMux
    port map (
            O => \N__21586\,
            I => \N__21564\
        );

    \I__2402\ : InMux
    port map (
            O => \N__21585\,
            I => \N__21564\
        );

    \I__2401\ : InMux
    port map (
            O => \N__21584\,
            I => \N__21561\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__21573\,
            I => \N__21558\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__21564\,
            I => \N__21555\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__21561\,
            I => \N__21548\
        );

    \I__2397\ : Span4Mux_v
    port map (
            O => \N__21558\,
            I => \N__21548\
        );

    \I__2396\ : Span4Mux_s3_h
    port map (
            O => \N__21555\,
            I => \N__21548\
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__21548\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2394\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21542\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__21542\,
            I => \N__21539\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__21539\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2391\ : CascadeMux
    port map (
            O => \N__21536\,
            I => \N__21533\
        );

    \I__2390\ : InMux
    port map (
            O => \N__21533\,
            I => \N__21530\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__21530\,
            I => \N__21527\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__21527\,
            I => \pwm_generator_inst.threshold_2\
        );

    \I__2387\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21521\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__21521\,
            I => \N__21517\
        );

    \I__2385\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21513\
        );

    \I__2384\ : Span4Mux_h
    port map (
            O => \N__21517\,
            I => \N__21510\
        );

    \I__2383\ : InMux
    port map (
            O => \N__21516\,
            I => \N__21507\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__21513\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__21510\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__21507\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2379\ : InMux
    port map (
            O => \N__21500\,
            I => \N__21497\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__21497\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2377\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21490\
        );

    \I__2376\ : InMux
    port map (
            O => \N__21493\,
            I => \N__21486\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__21490\,
            I => \N__21483\
        );

    \I__2374\ : InMux
    port map (
            O => \N__21489\,
            I => \N__21480\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__21486\,
            I => \N__21475\
        );

    \I__2372\ : Span4Mux_v
    port map (
            O => \N__21483\,
            I => \N__21475\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__21480\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2370\ : Odrv4
    port map (
            O => \N__21475\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__21470\,
            I => \N__21467\
        );

    \I__2368\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21464\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__21464\,
            I => \N__21461\
        );

    \I__2366\ : Odrv12
    port map (
            O => \N__21461\,
            I => \pwm_generator_inst.threshold_3\
        );

    \I__2365\ : InMux
    port map (
            O => \N__21458\,
            I => \N__21455\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__21455\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2363\ : InMux
    port map (
            O => \N__21452\,
            I => \N__21449\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__21449\,
            I => \N__21444\
        );

    \I__2361\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21441\
        );

    \I__2360\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21438\
        );

    \I__2359\ : Span4Mux_v
    port map (
            O => \N__21444\,
            I => \N__21435\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__21441\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__21438\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__21435\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2355\ : CascadeMux
    port map (
            O => \N__21428\,
            I => \N__21425\
        );

    \I__2354\ : InMux
    port map (
            O => \N__21425\,
            I => \N__21422\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__21422\,
            I => \pwm_generator_inst.threshold_4\
        );

    \I__2352\ : InMux
    port map (
            O => \N__21419\,
            I => \N__21416\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__21416\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__21413\,
            I => \N__21410\
        );

    \I__2349\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21407\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__21407\,
            I => \N__21404\
        );

    \I__2347\ : Odrv4
    port map (
            O => \N__21404\,
            I => \pwm_generator_inst.threshold_5\
        );

    \I__2346\ : InMux
    port map (
            O => \N__21401\,
            I => \N__21398\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__21398\,
            I => \N__21393\
        );

    \I__2344\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21390\
        );

    \I__2343\ : InMux
    port map (
            O => \N__21396\,
            I => \N__21387\
        );

    \I__2342\ : Span4Mux_v
    port map (
            O => \N__21393\,
            I => \N__21384\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__21390\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__21387\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__21384\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2338\ : InMux
    port map (
            O => \N__21377\,
            I => \N__21374\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__21374\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__21371\,
            I => \N__21368\
        );

    \I__2335\ : InMux
    port map (
            O => \N__21368\,
            I => \N__21365\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__21365\,
            I => \pwm_generator_inst.un14_counter_6\
        );

    \I__2333\ : InMux
    port map (
            O => \N__21362\,
            I => \N__21359\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__21359\,
            I => \N__21354\
        );

    \I__2331\ : InMux
    port map (
            O => \N__21358\,
            I => \N__21351\
        );

    \I__2330\ : InMux
    port map (
            O => \N__21357\,
            I => \N__21348\
        );

    \I__2329\ : Span4Mux_h
    port map (
            O => \N__21354\,
            I => \N__21345\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__21351\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__21348\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__21345\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2325\ : InMux
    port map (
            O => \N__21338\,
            I => \N__21335\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__21335\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__21332\,
            I => \N__21329\
        );

    \I__2322\ : InMux
    port map (
            O => \N__21329\,
            I => \N__21326\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__21326\,
            I => \pwm_generator_inst.un14_counter_7\
        );

    \I__2320\ : InMux
    port map (
            O => \N__21323\,
            I => \N__21320\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__21320\,
            I => \N__21315\
        );

    \I__2318\ : InMux
    port map (
            O => \N__21319\,
            I => \N__21312\
        );

    \I__2317\ : InMux
    port map (
            O => \N__21318\,
            I => \N__21309\
        );

    \I__2316\ : Span4Mux_v
    port map (
            O => \N__21315\,
            I => \N__21306\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__21312\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__21309\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2313\ : Odrv4
    port map (
            O => \N__21306\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2312\ : InMux
    port map (
            O => \N__21299\,
            I => \N__21296\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__21296\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__21293\,
            I => \N__21290\
        );

    \I__2309\ : InMux
    port map (
            O => \N__21290\,
            I => \N__21287\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__21287\,
            I => \pwm_generator_inst.un14_counter_8\
        );

    \I__2307\ : InMux
    port map (
            O => \N__21284\,
            I => \N__21281\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__21281\,
            I => \N__21277\
        );

    \I__2305\ : InMux
    port map (
            O => \N__21280\,
            I => \N__21273\
        );

    \I__2304\ : Span4Mux_h
    port map (
            O => \N__21277\,
            I => \N__21270\
        );

    \I__2303\ : InMux
    port map (
            O => \N__21276\,
            I => \N__21267\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__21273\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__21270\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__21267\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2299\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21257\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__21257\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__2296\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21248\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__21248\,
            I => \N__21245\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__21245\,
            I => \pwm_generator_inst.threshold_0\
        );

    \I__2293\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21239\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__21239\,
            I => \N__21235\
        );

    \I__2291\ : InMux
    port map (
            O => \N__21238\,
            I => \N__21231\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__21235\,
            I => \N__21228\
        );

    \I__2289\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21225\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__21231\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__21228\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__21225\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2285\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__21215\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__21212\,
            I => \N__21209\
        );

    \I__2282\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21206\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__21206\,
            I => \N__21203\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__21203\,
            I => \pwm_generator_inst.un14_counter_1\
        );

    \I__2279\ : InMux
    port map (
            O => \N__21200\,
            I => \N__21197\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__21197\,
            I => \N__21192\
        );

    \I__2277\ : InMux
    port map (
            O => \N__21196\,
            I => \N__21189\
        );

    \I__2276\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21186\
        );

    \I__2275\ : Span4Mux_h
    port map (
            O => \N__21192\,
            I => \N__21183\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__21189\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__21186\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__21183\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2271\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21172\
        );

    \I__2270\ : InMux
    port map (
            O => \N__21175\,
            I => \N__21169\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__21172\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__21169\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__2267\ : InMux
    port map (
            O => \N__21164\,
            I => \N__21161\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__21161\,
            I => \N__21156\
        );

    \I__2265\ : InMux
    port map (
            O => \N__21160\,
            I => \N__21151\
        );

    \I__2264\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21151\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__21156\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__21151\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__21146\,
            I => \N__21142\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__21145\,
            I => \N__21139\
        );

    \I__2259\ : InMux
    port map (
            O => \N__21142\,
            I => \N__21136\
        );

    \I__2258\ : InMux
    port map (
            O => \N__21139\,
            I => \N__21133\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__21136\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__21133\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__2255\ : InMux
    port map (
            O => \N__21128\,
            I => \N__21125\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__21125\,
            I => \N__21122\
        );

    \I__2253\ : Span4Mux_s2_h
    port map (
            O => \N__21122\,
            I => \N__21117\
        );

    \I__2252\ : InMux
    port map (
            O => \N__21121\,
            I => \N__21112\
        );

    \I__2251\ : InMux
    port map (
            O => \N__21120\,
            I => \N__21112\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__21117\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__21112\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2248\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21104\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__2246\ : Odrv12
    port map (
            O => \N__21101\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__2245\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21094\
        );

    \I__2244\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21091\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__21094\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__21091\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__2241\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21083\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__21083\,
            I => \N__21078\
        );

    \I__2239\ : InMux
    port map (
            O => \N__21082\,
            I => \N__21073\
        );

    \I__2238\ : InMux
    port map (
            O => \N__21081\,
            I => \N__21073\
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__21078\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__21073\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2235\ : InMux
    port map (
            O => \N__21068\,
            I => \N__21065\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__21065\,
            I => \N__21062\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__21062\,
            I => un7_start_stop
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__21059\,
            I => \N__21056\
        );

    \I__2231\ : InMux
    port map (
            O => \N__21056\,
            I => \N__21051\
        );

    \I__2230\ : InMux
    port map (
            O => \N__21055\,
            I => \N__21048\
        );

    \I__2229\ : InMux
    port map (
            O => \N__21054\,
            I => \N__21045\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__21051\,
            I => \N__21042\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__21048\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__21045\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__2225\ : Odrv12
    port map (
            O => \N__21042\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__2224\ : InMux
    port map (
            O => \N__21035\,
            I => \N__21032\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__21032\,
            I => \N__21029\
        );

    \I__2222\ : Span4Mux_s3_h
    port map (
            O => \N__21029\,
            I => \N__21026\
        );

    \I__2221\ : Odrv4
    port map (
            O => \N__21026\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\
        );

    \I__2220\ : InMux
    port map (
            O => \N__21023\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11\
        );

    \I__2219\ : InMux
    port map (
            O => \N__21020\,
            I => \N__21017\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__21017\,
            I => \N__21012\
        );

    \I__2217\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21009\
        );

    \I__2216\ : InMux
    port map (
            O => \N__21015\,
            I => \N__21006\
        );

    \I__2215\ : Sp12to4
    port map (
            O => \N__21012\,
            I => \N__21001\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__21009\,
            I => \N__21001\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__21006\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__2212\ : Odrv12
    port map (
            O => \N__21001\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__2211\ : InMux
    port map (
            O => \N__20996\,
            I => \N__20993\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__20993\,
            I => \N__20990\
        );

    \I__2209\ : Span4Mux_s3_h
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__2208\ : Odrv4
    port map (
            O => \N__20987\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\
        );

    \I__2207\ : InMux
    port map (
            O => \N__20984\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12\
        );

    \I__2206\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20978\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__20978\,
            I => \N__20973\
        );

    \I__2204\ : InMux
    port map (
            O => \N__20977\,
            I => \N__20970\
        );

    \I__2203\ : InMux
    port map (
            O => \N__20976\,
            I => \N__20967\
        );

    \I__2202\ : Span4Mux_v
    port map (
            O => \N__20973\,
            I => \N__20964\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__20970\,
            I => \N__20961\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__20967\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__20964\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__20961\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20954\,
            I => \N__20951\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__20951\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\
        );

    \I__2195\ : InMux
    port map (
            O => \N__20948\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__20945\,
            I => \N__20940\
        );

    \I__2193\ : InMux
    port map (
            O => \N__20944\,
            I => \N__20937\
        );

    \I__2192\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20934\
        );

    \I__2191\ : InMux
    port map (
            O => \N__20940\,
            I => \N__20931\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__20937\,
            I => \N__20928\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__20934\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__20931\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2187\ : Odrv4
    port map (
            O => \N__20928\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2186\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20918\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__20918\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\
        );

    \I__2184\ : InMux
    port map (
            O => \N__20915\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14\
        );

    \I__2183\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20909\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__20906\,
            I => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\
        );

    \I__2180\ : InMux
    port map (
            O => \N__20903\,
            I => \bfn_2_23_0_\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__20900\,
            I => \N__20897\
        );

    \I__2178\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20894\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__20894\,
            I => \N__20891\
        );

    \I__2176\ : Span4Mux_s2_h
    port map (
            O => \N__20891\,
            I => \N__20888\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__20888\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\
        );

    \I__2174\ : InMux
    port map (
            O => \N__20885\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16\
        );

    \I__2173\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__20879\,
            I => \N__20876\
        );

    \I__2171\ : Odrv4
    port map (
            O => \N__20876\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20873\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17\
        );

    \I__2169\ : InMux
    port map (
            O => \N__20870\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18\
        );

    \I__2168\ : InMux
    port map (
            O => \N__20867\,
            I => \N__20864\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__20864\,
            I => \N__20861\
        );

    \I__2166\ : Span4Mux_v
    port map (
            O => \N__20861\,
            I => \N__20858\
        );

    \I__2165\ : Odrv4
    port map (
            O => \N__20858\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\
        );

    \I__2164\ : InMux
    port map (
            O => \N__20855\,
            I => \N__20852\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__20852\,
            I => \N__20849\
        );

    \I__2162\ : Span4Mux_h
    port map (
            O => \N__20849\,
            I => \N__20846\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__20846\,
            I => \pwm_generator_inst.O_4\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20840\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__20840\,
            I => \pwm_generator_inst.un15_threshold_1_axb_4\
        );

    \I__2158\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20834\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__20834\,
            I => \N__20831\
        );

    \I__2156\ : Span4Mux_h
    port map (
            O => \N__20831\,
            I => \N__20828\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__20828\,
            I => \pwm_generator_inst.O_5\
        );

    \I__2154\ : InMux
    port map (
            O => \N__20825\,
            I => \N__20822\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__20822\,
            I => \pwm_generator_inst.un15_threshold_1_axb_5\
        );

    \I__2152\ : InMux
    port map (
            O => \N__20819\,
            I => \N__20816\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__20816\,
            I => \N__20813\
        );

    \I__2150\ : Span4Mux_h
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__20810\,
            I => \pwm_generator_inst.O_6\
        );

    \I__2148\ : InMux
    port map (
            O => \N__20807\,
            I => \N__20804\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__20804\,
            I => \pwm_generator_inst.un15_threshold_1_axb_6\
        );

    \I__2146\ : InMux
    port map (
            O => \N__20801\,
            I => \N__20798\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__20798\,
            I => \N__20795\
        );

    \I__2144\ : Span4Mux_h
    port map (
            O => \N__20795\,
            I => \N__20792\
        );

    \I__2143\ : Odrv4
    port map (
            O => \N__20792\,
            I => \pwm_generator_inst.O_7\
        );

    \I__2142\ : InMux
    port map (
            O => \N__20789\,
            I => \N__20786\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__20786\,
            I => \pwm_generator_inst.un15_threshold_1_axb_7\
        );

    \I__2140\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20780\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__2138\ : Span4Mux_h
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__20774\,
            I => \pwm_generator_inst.O_8\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20768\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__20768\,
            I => \pwm_generator_inst.un15_threshold_1_axb_8\
        );

    \I__2134\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20762\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__20762\,
            I => \N__20759\
        );

    \I__2132\ : Span4Mux_h
    port map (
            O => \N__20759\,
            I => \N__20756\
        );

    \I__2131\ : Odrv4
    port map (
            O => \N__20756\,
            I => \pwm_generator_inst.O_9\
        );

    \I__2130\ : InMux
    port map (
            O => \N__20753\,
            I => \N__20750\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__20750\,
            I => \pwm_generator_inst.un15_threshold_1_axb_9\
        );

    \I__2128\ : InMux
    port map (
            O => \N__20747\,
            I => \N__20742\
        );

    \I__2127\ : InMux
    port map (
            O => \N__20746\,
            I => \N__20739\
        );

    \I__2126\ : InMux
    port map (
            O => \N__20745\,
            I => \N__20736\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__20742\,
            I => \N__20733\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__20739\,
            I => \N__20730\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__20736\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__20733\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__2121\ : Odrv12
    port map (
            O => \N__20730\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__2120\ : InMux
    port map (
            O => \N__20723\,
            I => \N__20720\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__20720\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\
        );

    \I__2118\ : InMux
    port map (
            O => \N__20717\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9\
        );

    \I__2117\ : CascadeMux
    port map (
            O => \N__20714\,
            I => \N__20710\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__20713\,
            I => \N__20704\
        );

    \I__2115\ : InMux
    port map (
            O => \N__20710\,
            I => \N__20699\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__20709\,
            I => \N__20696\
        );

    \I__2113\ : CascadeMux
    port map (
            O => \N__20708\,
            I => \N__20692\
        );

    \I__2112\ : InMux
    port map (
            O => \N__20707\,
            I => \N__20686\
        );

    \I__2111\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20683\
        );

    \I__2110\ : InMux
    port map (
            O => \N__20703\,
            I => \N__20678\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20678\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__20699\,
            I => \N__20675\
        );

    \I__2107\ : InMux
    port map (
            O => \N__20696\,
            I => \N__20668\
        );

    \I__2106\ : InMux
    port map (
            O => \N__20695\,
            I => \N__20668\
        );

    \I__2105\ : InMux
    port map (
            O => \N__20692\,
            I => \N__20668\
        );

    \I__2104\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20665\
        );

    \I__2103\ : InMux
    port map (
            O => \N__20690\,
            I => \N__20660\
        );

    \I__2102\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20660\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__20686\,
            I => \N__20655\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__20683\,
            I => \N__20655\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__20678\,
            I => \N__20652\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__20675\,
            I => \N__20645\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__20668\,
            I => \N__20645\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__20665\,
            I => \N__20645\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__20660\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__2094\ : Odrv12
    port map (
            O => \N__20655\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__2093\ : Odrv4
    port map (
            O => \N__20652\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__20645\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__2091\ : InMux
    port map (
            O => \N__20636\,
            I => \N__20633\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__20633\,
            I => \N__20629\
        );

    \I__2089\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20626\
        );

    \I__2088\ : Span4Mux_v
    port map (
            O => \N__20629\,
            I => \N__20623\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__20626\,
            I => \N__20620\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__20623\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__20620\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__2084\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20612\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__20612\,
            I => \N__20609\
        );

    \I__2082\ : Span4Mux_v
    port map (
            O => \N__20609\,
            I => \N__20606\
        );

    \I__2081\ : Odrv4
    port map (
            O => \N__20606\,
            I => \pwm_generator_inst.un19_threshold_axb_1\
        );

    \I__2080\ : InMux
    port map (
            O => \N__20603\,
            I => \pwm_generator_inst.un15_threshold_1_cry_10\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__20600\,
            I => \N__20597\
        );

    \I__2078\ : InMux
    port map (
            O => \N__20597\,
            I => \N__20593\
        );

    \I__2077\ : InMux
    port map (
            O => \N__20596\,
            I => \N__20590\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__20593\,
            I => \N__20585\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__20590\,
            I => \N__20585\
        );

    \I__2074\ : Span4Mux_h
    port map (
            O => \N__20585\,
            I => \N__20582\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__20582\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__2072\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20575\
        );

    \I__2071\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20572\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__20575\,
            I => \N__20569\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__20572\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__20569\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__20564\,
            I => \N__20557\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__20563\,
            I => \N__20554\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__20562\,
            I => \N__20550\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__20561\,
            I => \N__20547\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__20560\,
            I => \N__20544\
        );

    \I__2062\ : InMux
    port map (
            O => \N__20557\,
            I => \N__20533\
        );

    \I__2061\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20533\
        );

    \I__2060\ : InMux
    port map (
            O => \N__20553\,
            I => \N__20533\
        );

    \I__2059\ : InMux
    port map (
            O => \N__20550\,
            I => \N__20533\
        );

    \I__2058\ : InMux
    port map (
            O => \N__20547\,
            I => \N__20533\
        );

    \I__2057\ : InMux
    port map (
            O => \N__20544\,
            I => \N__20526\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__20533\,
            I => \N__20523\
        );

    \I__2055\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20514\
        );

    \I__2054\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20514\
        );

    \I__2053\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20514\
        );

    \I__2052\ : InMux
    port map (
            O => \N__20529\,
            I => \N__20514\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__20526\,
            I => \N__20507\
        );

    \I__2050\ : Span4Mux_h
    port map (
            O => \N__20523\,
            I => \N__20507\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__20514\,
            I => \N__20507\
        );

    \I__2048\ : Odrv4
    port map (
            O => \N__20507\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2047\ : InMux
    port map (
            O => \N__20504\,
            I => \N__20500\
        );

    \I__2046\ : InMux
    port map (
            O => \N__20503\,
            I => \N__20497\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__20500\,
            I => \N__20494\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__20497\,
            I => \N__20491\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__20494\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__20491\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__2041\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20483\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__20483\,
            I => \N__20480\
        );

    \I__2039\ : Span4Mux_v
    port map (
            O => \N__20480\,
            I => \N__20477\
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__20477\,
            I => \pwm_generator_inst.O_0\
        );

    \I__2037\ : InMux
    port map (
            O => \N__20474\,
            I => \N__20471\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__20471\,
            I => \pwm_generator_inst.un15_threshold_1_axb_0\
        );

    \I__2035\ : InMux
    port map (
            O => \N__20468\,
            I => \N__20465\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__20465\,
            I => \N__20462\
        );

    \I__2033\ : Span4Mux_h
    port map (
            O => \N__20462\,
            I => \N__20459\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__20459\,
            I => \pwm_generator_inst.O_1\
        );

    \I__2031\ : InMux
    port map (
            O => \N__20456\,
            I => \N__20453\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__20453\,
            I => \pwm_generator_inst.un15_threshold_1_axb_1\
        );

    \I__2029\ : InMux
    port map (
            O => \N__20450\,
            I => \N__20447\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__20447\,
            I => \N__20444\
        );

    \I__2027\ : Span4Mux_v
    port map (
            O => \N__20444\,
            I => \N__20441\
        );

    \I__2026\ : Odrv4
    port map (
            O => \N__20441\,
            I => \pwm_generator_inst.O_2\
        );

    \I__2025\ : InMux
    port map (
            O => \N__20438\,
            I => \N__20435\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__20435\,
            I => \pwm_generator_inst.un15_threshold_1_axb_2\
        );

    \I__2023\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20429\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__20429\,
            I => \N__20426\
        );

    \I__2021\ : Span4Mux_v
    port map (
            O => \N__20426\,
            I => \N__20423\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__20423\,
            I => \pwm_generator_inst.O_3\
        );

    \I__2019\ : InMux
    port map (
            O => \N__20420\,
            I => \N__20417\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__20417\,
            I => \pwm_generator_inst.un15_threshold_1_axb_3\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__2016\ : InMux
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__20408\,
            I => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\
        );

    \I__2014\ : InMux
    port map (
            O => \N__20405\,
            I => \N__20402\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__20402\,
            I => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\
        );

    \I__2012\ : InMux
    port map (
            O => \N__20399\,
            I => \N__20396\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__20396\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__2009\ : InMux
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__20387\,
            I => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\
        );

    \I__2007\ : InMux
    port map (
            O => \N__20384\,
            I => \N__20381\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__20381\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\
        );

    \I__2005\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20375\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__20375\,
            I => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\
        );

    \I__2003\ : InMux
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__20369\,
            I => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__20366\,
            I => \N__20358\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__20365\,
            I => \N__20354\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__20364\,
            I => \N__20351\
        );

    \I__1998\ : InMux
    port map (
            O => \N__20363\,
            I => \N__20346\
        );

    \I__1997\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20346\
        );

    \I__1996\ : InMux
    port map (
            O => \N__20361\,
            I => \N__20340\
        );

    \I__1995\ : InMux
    port map (
            O => \N__20358\,
            I => \N__20310\
        );

    \I__1994\ : InMux
    port map (
            O => \N__20357\,
            I => \N__20310\
        );

    \I__1993\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20310\
        );

    \I__1992\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20310\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__20346\,
            I => \N__20307\
        );

    \I__1990\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20300\
        );

    \I__1989\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20300\
        );

    \I__1988\ : InMux
    port map (
            O => \N__20343\,
            I => \N__20300\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__20340\,
            I => \N__20297\
        );

    \I__1986\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20286\
        );

    \I__1985\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20286\
        );

    \I__1984\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20286\
        );

    \I__1983\ : InMux
    port map (
            O => \N__20336\,
            I => \N__20286\
        );

    \I__1982\ : InMux
    port map (
            O => \N__20335\,
            I => \N__20286\
        );

    \I__1981\ : InMux
    port map (
            O => \N__20334\,
            I => \N__20268\
        );

    \I__1980\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20268\
        );

    \I__1979\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20268\
        );

    \I__1978\ : InMux
    port map (
            O => \N__20331\,
            I => \N__20268\
        );

    \I__1977\ : InMux
    port map (
            O => \N__20330\,
            I => \N__20268\
        );

    \I__1976\ : InMux
    port map (
            O => \N__20329\,
            I => \N__20268\
        );

    \I__1975\ : InMux
    port map (
            O => \N__20328\,
            I => \N__20268\
        );

    \I__1974\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20268\
        );

    \I__1973\ : InMux
    port map (
            O => \N__20326\,
            I => \N__20253\
        );

    \I__1972\ : InMux
    port map (
            O => \N__20325\,
            I => \N__20253\
        );

    \I__1971\ : InMux
    port map (
            O => \N__20324\,
            I => \N__20253\
        );

    \I__1970\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20253\
        );

    \I__1969\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20253\
        );

    \I__1968\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20253\
        );

    \I__1967\ : InMux
    port map (
            O => \N__20320\,
            I => \N__20253\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__20319\,
            I => \N__20250\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__20310\,
            I => \N__20247\
        );

    \I__1964\ : Span4Mux_s1_h
    port map (
            O => \N__20307\,
            I => \N__20242\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__20300\,
            I => \N__20242\
        );

    \I__1962\ : Span4Mux_v
    port map (
            O => \N__20297\,
            I => \N__20237\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__20286\,
            I => \N__20237\
        );

    \I__1960\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20234\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__20268\,
            I => \N__20229\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__20253\,
            I => \N__20229\
        );

    \I__1957\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20226\
        );

    \I__1956\ : Span4Mux_h
    port map (
            O => \N__20247\,
            I => \N__20221\
        );

    \I__1955\ : Span4Mux_v
    port map (
            O => \N__20242\,
            I => \N__20221\
        );

    \I__1954\ : Span4Mux_v
    port map (
            O => \N__20237\,
            I => \N__20218\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__20234\,
            I => \N__20215\
        );

    \I__1952\ : Span4Mux_s1_h
    port map (
            O => \N__20229\,
            I => \N__20212\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__20226\,
            I => \N__20207\
        );

    \I__1950\ : Sp12to4
    port map (
            O => \N__20221\,
            I => \N__20207\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__20218\,
            I => \N_19_1\
        );

    \I__1948\ : Odrv12
    port map (
            O => \N__20215\,
            I => \N_19_1\
        );

    \I__1947\ : Odrv4
    port map (
            O => \N__20212\,
            I => \N_19_1\
        );

    \I__1946\ : Odrv12
    port map (
            O => \N__20207\,
            I => \N_19_1\
        );

    \I__1945\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20195\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__20195\,
            I => \N__20191\
        );

    \I__1943\ : InMux
    port map (
            O => \N__20194\,
            I => \N__20188\
        );

    \I__1942\ : Span4Mux_v
    port map (
            O => \N__20191\,
            I => \N__20185\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__20188\,
            I => \N__20182\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__20185\,
            I => \N__20179\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__20182\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__20179\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__20174\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__20171\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__1935\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20150\
        );

    \I__1934\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20150\
        );

    \I__1933\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20150\
        );

    \I__1932\ : InMux
    port map (
            O => \N__20165\,
            I => \N__20150\
        );

    \I__1931\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20145\
        );

    \I__1930\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20145\
        );

    \I__1929\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20136\
        );

    \I__1928\ : InMux
    port map (
            O => \N__20161\,
            I => \N__20136\
        );

    \I__1927\ : InMux
    port map (
            O => \N__20160\,
            I => \N__20136\
        );

    \I__1926\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20136\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__20150\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__20145\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__20136\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__1922\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20126\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__20126\,
            I => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__20123\,
            I => \N__20120\
        );

    \I__1919\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20116\
        );

    \I__1918\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20113\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__20116\,
            I => \N__20108\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__20113\,
            I => \N__20108\
        );

    \I__1915\ : Span4Mux_v
    port map (
            O => \N__20108\,
            I => \N__20105\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__20105\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__1913\ : InMux
    port map (
            O => \N__20102\,
            I => \N__20099\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__20099\,
            I => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\
        );

    \I__1911\ : InMux
    port map (
            O => \N__20096\,
            I => \N__20093\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__20093\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__1909\ : InMux
    port map (
            O => \N__20090\,
            I => \N__20087\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__20087\,
            I => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\
        );

    \I__1907\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20081\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__1905\ : Odrv12
    port map (
            O => \N__20078\,
            I => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\
        );

    \I__1904\ : InMux
    port map (
            O => \N__20075\,
            I => \N__20072\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__20072\,
            I => \N__20069\
        );

    \I__1902\ : Odrv12
    port map (
            O => \N__20069\,
            I => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\
        );

    \I__1901\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20063\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__20063\,
            I => \N__20060\
        );

    \I__1899\ : Odrv12
    port map (
            O => \N__20060\,
            I => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\
        );

    \I__1898\ : InMux
    port map (
            O => \N__20057\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__1897\ : InMux
    port map (
            O => \N__20054\,
            I => \N__20051\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__20051\,
            I => \N__20048\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__20048\,
            I => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\
        );

    \I__1894\ : InMux
    port map (
            O => \N__20045\,
            I => \N__20042\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__20042\,
            I => \N_86_i_i\
        );

    \I__1892\ : InMux
    port map (
            O => \N__20039\,
            I => \bfn_1_23_0_\
        );

    \I__1891\ : InMux
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__20027\,
            I => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\
        );

    \I__1887\ : InMux
    port map (
            O => \N__20024\,
            I => \N__20021\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__20021\,
            I => \N__20018\
        );

    \I__1885\ : Odrv12
    port map (
            O => \N__20018\,
            I => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\
        );

    \I__1884\ : InMux
    port map (
            O => \N__20015\,
            I => \N__20012\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__20012\,
            I => \N__20009\
        );

    \I__1882\ : Odrv12
    port map (
            O => \N__20009\,
            I => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\
        );

    \I__1881\ : InMux
    port map (
            O => \N__20006\,
            I => \N__20003\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__20003\,
            I => \N__20000\
        );

    \I__1879\ : Odrv12
    port map (
            O => \N__20000\,
            I => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\
        );

    \I__1878\ : InMux
    port map (
            O => \N__19997\,
            I => \N__19994\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__19994\,
            I => \N__19991\
        );

    \I__1876\ : Odrv12
    port map (
            O => \N__19991\,
            I => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\
        );

    \I__1875\ : InMux
    port map (
            O => \N__19988\,
            I => \N__19985\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__1873\ : Odrv4
    port map (
            O => \N__19982\,
            I => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\
        );

    \I__1872\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19976\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__19976\,
            I => \N__19973\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__19973\,
            I => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\
        );

    \I__1869\ : InMux
    port map (
            O => \N__19970\,
            I => \N__19967\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__19967\,
            I => \N__19964\
        );

    \I__1867\ : Odrv12
    port map (
            O => \N__19964\,
            I => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\
        );

    \I__1866\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__19958\,
            I => \N__19955\
        );

    \I__1864\ : Odrv4
    port map (
            O => \N__19955\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1863\ : InMux
    port map (
            O => \N__19952\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__1862\ : InMux
    port map (
            O => \N__19949\,
            I => \N__19946\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__19946\,
            I => \N__19943\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__19943\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1859\ : InMux
    port map (
            O => \N__19940\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__1858\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__19931\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1855\ : InMux
    port map (
            O => \N__19928\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__1854\ : InMux
    port map (
            O => \N__19925\,
            I => \N__19922\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__1852\ : Span4Mux_v
    port map (
            O => \N__19919\,
            I => \N__19916\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__19916\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_4\
        );

    \I__1850\ : InMux
    port map (
            O => \N__19913\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__19910\,
            I => \N__19907\
        );

    \I__1848\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19904\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__19904\,
            I => \N__19901\
        );

    \I__1846\ : Odrv12
    port map (
            O => \N__19901\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\
        );

    \I__1845\ : InMux
    port map (
            O => \N__19898\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__1844\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__19889\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\
        );

    \I__1841\ : InMux
    port map (
            O => \N__19886\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__19883\,
            I => \N__19880\
        );

    \I__1839\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__1837\ : Odrv4
    port map (
            O => \N__19874\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\
        );

    \I__1836\ : InMux
    port map (
            O => \N__19871\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__1835\ : InMux
    port map (
            O => \N__19868\,
            I => \N__19865\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__19865\,
            I => \N__19862\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__19862\,
            I => \N__19859\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__19859\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\
        );

    \I__1831\ : InMux
    port map (
            O => \N__19856\,
            I => \N__19853\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__1829\ : Span4Mux_v
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__1828\ : Odrv4
    port map (
            O => \N__19847\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\
        );

    \I__1827\ : InMux
    port map (
            O => \N__19844\,
            I => \N__19841\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__19841\,
            I => \N__19838\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__19838\,
            I => \N__19835\
        );

    \I__1824\ : Span4Mux_v
    port map (
            O => \N__19835\,
            I => \N__19832\
        );

    \I__1823\ : Span4Mux_v
    port map (
            O => \N__19832\,
            I => \N__19829\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__19829\,
            I => \pwm_generator_inst.un2_threshold_2_14\
        );

    \I__1821\ : InMux
    port map (
            O => \N__19826\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13\
        );

    \I__1820\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19820\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__19817\,
            I => \N__19813\
        );

    \I__1817\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19810\
        );

    \I__1816\ : Span4Mux_v
    port map (
            O => \N__19813\,
            I => \N__19802\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__19810\,
            I => \N__19802\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__19809\,
            I => \N__19798\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__19808\,
            I => \N__19794\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__19807\,
            I => \N__19790\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__19802\,
            I => \N__19787\
        );

    \I__1810\ : InMux
    port map (
            O => \N__19801\,
            I => \N__19774\
        );

    \I__1809\ : InMux
    port map (
            O => \N__19798\,
            I => \N__19774\
        );

    \I__1808\ : InMux
    port map (
            O => \N__19797\,
            I => \N__19774\
        );

    \I__1807\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19774\
        );

    \I__1806\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19774\
        );

    \I__1805\ : InMux
    port map (
            O => \N__19790\,
            I => \N__19774\
        );

    \I__1804\ : Span4Mux_v
    port map (
            O => \N__19787\,
            I => \N__19769\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__19774\,
            I => \N__19769\
        );

    \I__1802\ : Span4Mux_v
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__19766\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__1799\ : InMux
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__1797\ : Span12Mux_v
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__1796\ : Odrv12
    port map (
            O => \N__19751\,
            I => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\
        );

    \I__1795\ : InMux
    port map (
            O => \N__19748\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14\
        );

    \I__1794\ : InMux
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__19742\,
            I => \N__19739\
        );

    \I__1792\ : Odrv12
    port map (
            O => \N__19739\,
            I => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\
        );

    \I__1791\ : InMux
    port map (
            O => \N__19736\,
            I => \bfn_1_21_0_\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__19733\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81_cascade_\
        );

    \I__1789\ : InMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__19724\,
            I => \N__19721\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__19721\,
            I => \pwm_generator_inst.un19_threshold_axb_0\
        );

    \I__1785\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__1783\ : Odrv12
    port map (
            O => \N__19712\,
            I => \pwm_generator_inst.un19_threshold_axb_4\
        );

    \I__1782\ : InMux
    port map (
            O => \N__19709\,
            I => \N__19706\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__1780\ : Odrv12
    port map (
            O => \N__19703\,
            I => \pwm_generator_inst.un19_threshold_axb_5\
        );

    \I__1779\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19697\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__19697\,
            I => \N__19694\
        );

    \I__1777\ : Span4Mux_s2_h
    port map (
            O => \N__19694\,
            I => \N__19691\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__19691\,
            I => \pwm_generator_inst.un19_threshold_axb_6\
        );

    \I__1775\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19685\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__19685\,
            I => \N__19682\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__19682\,
            I => \pwm_generator_inst.un19_threshold_axb_8\
        );

    \I__1772\ : InMux
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__1770\ : Odrv12
    port map (
            O => \N__19673\,
            I => \pwm_generator_inst.un19_threshold_axb_7\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__19667\,
            I => \N__19664\
        );

    \I__1767\ : Span4Mux_v
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__1766\ : Span4Mux_v
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__1765\ : Span4Mux_v
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__19655\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__1763\ : CascadeMux
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__1762\ : InMux
    port map (
            O => \N__19649\,
            I => \N__19646\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__1760\ : Span4Mux_v
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__1759\ : Odrv4
    port map (
            O => \N__19640\,
            I => \pwm_generator_inst.un2_threshold_1_21\
        );

    \I__1758\ : InMux
    port map (
            O => \N__19637\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__1757\ : InMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__19631\,
            I => \N__19628\
        );

    \I__1755\ : Span4Mux_v
    port map (
            O => \N__19628\,
            I => \N__19625\
        );

    \I__1754\ : Span4Mux_v
    port map (
            O => \N__19625\,
            I => \N__19622\
        );

    \I__1753\ : Span4Mux_v
    port map (
            O => \N__19622\,
            I => \N__19619\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__19619\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__19616\,
            I => \N__19613\
        );

    \I__1750\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__19607\,
            I => \N__19604\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__19604\,
            I => \pwm_generator_inst.un2_threshold_1_22\
        );

    \I__1746\ : InMux
    port map (
            O => \N__19601\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__1745\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__1743\ : Span4Mux_v
    port map (
            O => \N__19592\,
            I => \N__19589\
        );

    \I__1742\ : Span4Mux_v
    port map (
            O => \N__19589\,
            I => \N__19586\
        );

    \I__1741\ : Span4Mux_v
    port map (
            O => \N__19586\,
            I => \N__19583\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__19583\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__1738\ : InMux
    port map (
            O => \N__19577\,
            I => \N__19574\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__19574\,
            I => \N__19571\
        );

    \I__1736\ : Span4Mux_v
    port map (
            O => \N__19571\,
            I => \N__19568\
        );

    \I__1735\ : Odrv4
    port map (
            O => \N__19568\,
            I => \pwm_generator_inst.un2_threshold_1_23\
        );

    \I__1734\ : InMux
    port map (
            O => \N__19565\,
            I => \bfn_1_20_0_\
        );

    \I__1733\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__19559\,
            I => \N__19556\
        );

    \I__1731\ : Span4Mux_v
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__1730\ : Span4Mux_v
    port map (
            O => \N__19553\,
            I => \N__19550\
        );

    \I__1729\ : Span4Mux_v
    port map (
            O => \N__19550\,
            I => \N__19547\
        );

    \I__1728\ : Odrv4
    port map (
            O => \N__19547\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__19544\,
            I => \N__19541\
        );

    \I__1726\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19538\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__1724\ : Span4Mux_v
    port map (
            O => \N__19535\,
            I => \N__19532\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__19532\,
            I => \pwm_generator_inst.un2_threshold_1_24\
        );

    \I__1722\ : InMux
    port map (
            O => \N__19529\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__1721\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__19523\,
            I => \N__19520\
        );

    \I__1719\ : Span12Mux_h
    port map (
            O => \N__19520\,
            I => \N__19517\
        );

    \I__1718\ : Span12Mux_v
    port map (
            O => \N__19517\,
            I => \N__19514\
        );

    \I__1717\ : Odrv12
    port map (
            O => \N__19514\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__1716\ : InMux
    port map (
            O => \N__19511\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__1715\ : CascadeMux
    port map (
            O => \N__19508\,
            I => \N__19505\
        );

    \I__1714\ : InMux
    port map (
            O => \N__19505\,
            I => \N__19502\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__19502\,
            I => \N__19499\
        );

    \I__1712\ : Span4Mux_h
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__19496\,
            I => \N__19493\
        );

    \I__1710\ : Sp12to4
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__1709\ : Odrv12
    port map (
            O => \N__19490\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__1708\ : InMux
    port map (
            O => \N__19487\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__1707\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19481\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__1705\ : Span4Mux_v
    port map (
            O => \N__19478\,
            I => \N__19475\
        );

    \I__1704\ : Span4Mux_v
    port map (
            O => \N__19475\,
            I => \N__19472\
        );

    \I__1703\ : Span4Mux_v
    port map (
            O => \N__19472\,
            I => \N__19469\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__19469\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__1701\ : InMux
    port map (
            O => \N__19466\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__1699\ : InMux
    port map (
            O => \N__19460\,
            I => \N__19457\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__19457\,
            I => \N__19454\
        );

    \I__1697\ : Span4Mux_h
    port map (
            O => \N__19454\,
            I => \N__19451\
        );

    \I__1696\ : Sp12to4
    port map (
            O => \N__19451\,
            I => \N__19448\
        );

    \I__1695\ : Span12Mux_v
    port map (
            O => \N__19448\,
            I => \N__19445\
        );

    \I__1694\ : Odrv12
    port map (
            O => \N__19445\,
            I => \pwm_generator_inst.un2_threshold_2_13\
        );

    \I__1693\ : InMux
    port map (
            O => \N__19442\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12\
        );

    \I__1692\ : InMux
    port map (
            O => \N__19439\,
            I => \N__19436\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__19436\,
            I => \pwm_generator_inst.un19_threshold_axb_2\
        );

    \I__1690\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19430\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__19430\,
            I => \pwm_generator_inst.un19_threshold_axb_3\
        );

    \I__1688\ : InMux
    port map (
            O => \N__19427\,
            I => \N__19424\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__19424\,
            I => \N__19421\
        );

    \I__1686\ : Span4Mux_v
    port map (
            O => \N__19421\,
            I => \N__19418\
        );

    \I__1685\ : Span4Mux_v
    port map (
            O => \N__19418\,
            I => \N__19415\
        );

    \I__1684\ : Span4Mux_v
    port map (
            O => \N__19415\,
            I => \N__19412\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__19412\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__19409\,
            I => \N__19406\
        );

    \I__1681\ : InMux
    port map (
            O => \N__19406\,
            I => \N__19403\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__19403\,
            I => \N__19400\
        );

    \I__1679\ : Span4Mux_v
    port map (
            O => \N__19400\,
            I => \N__19397\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__19397\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__1677\ : InMux
    port map (
            O => \N__19394\,
            I => \N__19391\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__19391\,
            I => \N__19388\
        );

    \I__1675\ : Span4Mux_v
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__1674\ : Span4Mux_v
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__1673\ : Span4Mux_v
    port map (
            O => \N__19382\,
            I => \N__19379\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__19379\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__1670\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__19370\,
            I => \N__19367\
        );

    \I__1668\ : Span4Mux_v
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__19364\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__1666\ : InMux
    port map (
            O => \N__19361\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__1665\ : InMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__19355\,
            I => \N__19352\
        );

    \I__1663\ : Span12Mux_h
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__1662\ : Span12Mux_v
    port map (
            O => \N__19349\,
            I => \N__19346\
        );

    \I__1661\ : Odrv12
    port map (
            O => \N__19346\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__19343\,
            I => \N__19340\
        );

    \I__1659\ : InMux
    port map (
            O => \N__19340\,
            I => \N__19337\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__19337\,
            I => \N__19334\
        );

    \I__1657\ : Span4Mux_v
    port map (
            O => \N__19334\,
            I => \N__19331\
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__19331\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__1655\ : InMux
    port map (
            O => \N__19328\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__1654\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19322\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__19322\,
            I => \N__19319\
        );

    \I__1652\ : Span4Mux_v
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__1651\ : Span4Mux_v
    port map (
            O => \N__19316\,
            I => \N__19313\
        );

    \I__1650\ : Span4Mux_v
    port map (
            O => \N__19313\,
            I => \N__19310\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__19310\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__19307\,
            I => \N__19304\
        );

    \I__1647\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__19301\,
            I => \N__19298\
        );

    \I__1645\ : Span4Mux_v
    port map (
            O => \N__19298\,
            I => \N__19295\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__19295\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__1643\ : InMux
    port map (
            O => \N__19292\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__1642\ : InMux
    port map (
            O => \N__19289\,
            I => \N__19286\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__19286\,
            I => \N__19283\
        );

    \I__1640\ : Span4Mux_v
    port map (
            O => \N__19283\,
            I => \N__19280\
        );

    \I__1639\ : Span4Mux_v
    port map (
            O => \N__19280\,
            I => \N__19277\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__19274\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__1635\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__19265\,
            I => \N__19262\
        );

    \I__1633\ : Span4Mux_v
    port map (
            O => \N__19262\,
            I => \N__19259\
        );

    \I__1632\ : Span4Mux_v
    port map (
            O => \N__19259\,
            I => \N__19256\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__19256\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__1630\ : InMux
    port map (
            O => \N__19253\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__1629\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19247\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__19247\,
            I => \N__19244\
        );

    \I__1627\ : Span4Mux_v
    port map (
            O => \N__19244\,
            I => \N__19241\
        );

    \I__1626\ : Span4Mux_v
    port map (
            O => \N__19241\,
            I => \N__19238\
        );

    \I__1625\ : Span4Mux_v
    port map (
            O => \N__19238\,
            I => \N__19235\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__19235\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__1622\ : InMux
    port map (
            O => \N__19229\,
            I => \N__19226\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__19226\,
            I => \N__19223\
        );

    \I__1620\ : Span4Mux_h
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__1619\ : Span4Mux_v
    port map (
            O => \N__19220\,
            I => \N__19217\
        );

    \I__1618\ : Odrv4
    port map (
            O => \N__19217\,
            I => \pwm_generator_inst.un2_threshold_1_20\
        );

    \I__1617\ : InMux
    port map (
            O => \N__19214\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__1616\ : InMux
    port map (
            O => \N__19211\,
            I => \pwm_generator_inst.un19_threshold_cry_0\
        );

    \I__1615\ : InMux
    port map (
            O => \N__19208\,
            I => \pwm_generator_inst.un19_threshold_cry_1\
        );

    \I__1614\ : InMux
    port map (
            O => \N__19205\,
            I => \pwm_generator_inst.un19_threshold_cry_2\
        );

    \I__1613\ : InMux
    port map (
            O => \N__19202\,
            I => \pwm_generator_inst.un19_threshold_cry_3\
        );

    \I__1612\ : InMux
    port map (
            O => \N__19199\,
            I => \pwm_generator_inst.un19_threshold_cry_4\
        );

    \I__1611\ : InMux
    port map (
            O => \N__19196\,
            I => \pwm_generator_inst.un19_threshold_cry_5\
        );

    \I__1610\ : InMux
    port map (
            O => \N__19193\,
            I => \pwm_generator_inst.un19_threshold_cry_6\
        );

    \I__1609\ : InMux
    port map (
            O => \N__19190\,
            I => \bfn_1_18_0_\
        );

    \I__1608\ : InMux
    port map (
            O => \N__19187\,
            I => \pwm_generator_inst.un19_threshold_cry_8\
        );

    \I__1607\ : InMux
    port map (
            O => \N__19184\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__1606\ : InMux
    port map (
            O => \N__19181\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__1605\ : InMux
    port map (
            O => \N__19178\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__1604\ : InMux
    port map (
            O => \N__19175\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__1603\ : InMux
    port map (
            O => \N__19172\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__1602\ : InMux
    port map (
            O => \N__19169\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__1601\ : InMux
    port map (
            O => \N__19166\,
            I => \bfn_1_16_0_\
        );

    \I__1600\ : InMux
    port map (
            O => \N__19163\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__1599\ : InMux
    port map (
            O => \N__19160\,
            I => \N__19157\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__19157\,
            I => \N__19154\
        );

    \I__1597\ : Span4Mux_v
    port map (
            O => \N__19154\,
            I => \N__19150\
        );

    \I__1596\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19147\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__19150\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__19147\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__1593\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19139\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__1591\ : Span4Mux_v
    port map (
            O => \N__19136\,
            I => \N__19133\
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__19133\,
            I => \pwm_generator_inst.un2_threshold_2_1_16\
        );

    \I__1589\ : InMux
    port map (
            O => \N__19130\,
            I => \bfn_1_15_0_\
        );

    \I__1588\ : InMux
    port map (
            O => \N__19127\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__1587\ : IoInMux
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__19121\,
            I => \N__19118\
        );

    \I__1585\ : Span4Mux_s3_v
    port map (
            O => \N__19118\,
            I => \N__19115\
        );

    \I__1584\ : Span4Mux_h
    port map (
            O => \N__19115\,
            I => \N__19112\
        );

    \I__1583\ : Sp12to4
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__1582\ : Span12Mux_v
    port map (
            O => \N__19109\,
            I => \N__19106\
        );

    \I__1581\ : Span12Mux_v
    port map (
            O => \N__19106\,
            I => \N__19103\
        );

    \I__1580\ : Odrv12
    port map (
            O => \N__19103\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1579\ : IoInMux
    port map (
            O => \N__19100\,
            I => \N__19097\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__19097\,
            I => \N__19094\
        );

    \I__1577\ : IoSpan4Mux
    port map (
            O => \N__19094\,
            I => \N__19091\
        );

    \I__1576\ : IoSpan4Mux
    port map (
            O => \N__19091\,
            I => \N__19088\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__19088\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_1_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_22_0_\
        );

    \IN_MUX_bfv_1_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_1_23_0_\
        );

    \IN_MUX_bfv_1_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_1_24_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_15_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_5_0_\
        );

    \IN_MUX_bfv_15_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_15_6_0_\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_4_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryinitout => \bfn_4_15_0_\
        );

    \IN_MUX_bfv_5_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_19_0_\
        );

    \IN_MUX_bfv_5_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryinitout => \bfn_5_20_0_\
        );

    \IN_MUX_bfv_5_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryinitout => \bfn_5_21_0_\
        );

    \IN_MUX_bfv_5_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryinitout => \bfn_5_22_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_1_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_1_20_0_\
        );

    \IN_MUX_bfv_1_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            carryinitout => \bfn_1_21_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_cry_7\,
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_2_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_21_0_\
        );

    \IN_MUX_bfv_2_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_7\,
            carryinitout => \bfn_2_22_0_\
        );

    \IN_MUX_bfv_2_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_15\,
            carryinitout => \bfn_2_23_0_\
        );

    \IN_MUX_bfv_3_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_16_0_\
        );

    \IN_MUX_bfv_3_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_3_17_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_15_12_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_10_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_10_11_0_\
        );

    \IN_MUX_bfv_14_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_4_0_\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_18_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_7_0_\
        );

    \IN_MUX_bfv_18_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_18_8_0_\
        );

    \IN_MUX_bfv_18_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_18_9_0_\
        );

    \IN_MUX_bfv_18_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_18_10_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_15\,
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_23\,
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_18_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_18_21_0_\
        );

    \IN_MUX_bfv_18_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_18_22_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_16_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_16_18_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_16_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_16_20_0_\
        );

    \IN_MUX_bfv_18_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_23_0_\
        );

    \IN_MUX_bfv_18_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_18_24_0_\
        );

    \IN_MUX_bfv_18_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_18_25_0_\
        );

    \IN_MUX_bfv_18_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_18_26_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_11_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            carryinitout => \bfn_11_21_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            carryinitout => \bfn_11_22_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19124\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19100\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__35834\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_161_i_g\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__26210\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__36881\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__44747\,
            CLKHFEN => \N__44786\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__44785\,
            RGB2PWM => \N__20045\,
            RGB1 => rgb_g_wire,
            CURREN => \N__44831\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__21068\,
            RGB0PWM => \N__49271\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__19823\,
            in1 => \N__19153\,
            in2 => \_gnd_net_\,
            in3 => \N__20285\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25250\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50049\,
            ce => 'H',
            sr => \N__49207\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__19160\,
            in1 => \N__19816\,
            in2 => \N__20319\,
            in3 => \N__19142\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20165\,
            in1 => \N__21238\,
            in2 => \_gnd_net_\,
            in3 => \N__19130\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__50020\,
            ce => 'H',
            sr => \N__49227\
        );

    \pwm_generator_inst.counter_1_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20159\,
            in1 => \N__21196\,
            in2 => \_gnd_net_\,
            in3 => \N__19127\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__50020\,
            ce => 'H',
            sr => \N__49227\
        );

    \pwm_generator_inst.counter_2_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20166\,
            in1 => \N__21520\,
            in2 => \_gnd_net_\,
            in3 => \N__19184\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__50020\,
            ce => 'H',
            sr => \N__49227\
        );

    \pwm_generator_inst.counter_3_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20160\,
            in1 => \N__21493\,
            in2 => \_gnd_net_\,
            in3 => \N__19181\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__50020\,
            ce => 'H',
            sr => \N__49227\
        );

    \pwm_generator_inst.counter_4_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20167\,
            in1 => \N__21448\,
            in2 => \_gnd_net_\,
            in3 => \N__19178\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__50020\,
            ce => 'H',
            sr => \N__49227\
        );

    \pwm_generator_inst.counter_5_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20161\,
            in1 => \N__21396\,
            in2 => \_gnd_net_\,
            in3 => \N__19175\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__50020\,
            ce => 'H',
            sr => \N__49227\
        );

    \pwm_generator_inst.counter_6_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20168\,
            in1 => \N__21357\,
            in2 => \_gnd_net_\,
            in3 => \N__19172\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__50020\,
            ce => 'H',
            sr => \N__49227\
        );

    \pwm_generator_inst.counter_7_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20162\,
            in1 => \N__21319\,
            in2 => \_gnd_net_\,
            in3 => \N__19169\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__50020\,
            ce => 'H',
            sr => \N__49227\
        );

    \pwm_generator_inst.counter_8_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20164\,
            in1 => \N__21280\,
            in2 => \_gnd_net_\,
            in3 => \N__19166\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__50010\,
            ce => 'H',
            sr => \N__49233\
        );

    \pwm_generator_inst.counter_9_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21649\,
            in1 => \N__20163\,
            in2 => \_gnd_net_\,
            in3 => \N__19163\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50010\,
            ce => 'H',
            sr => \N__49233\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19730\,
            in2 => \N__20713\,
            in3 => \N__20707\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20615\,
            in2 => \_gnd_net_\,
            in3 => \N__19211\,
            lcout => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19439\,
            in2 => \_gnd_net_\,
            in3 => \N__19208\,
            lcout => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19433\,
            in2 => \_gnd_net_\,
            in3 => \N__19205\,
            lcout => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19718\,
            in2 => \_gnd_net_\,
            in3 => \N__19202\,
            lcout => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19709\,
            in2 => \_gnd_net_\,
            in3 => \N__19199\,
            lcout => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19700\,
            in2 => \_gnd_net_\,
            in3 => \N__19196\,
            lcout => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19679\,
            in2 => \_gnd_net_\,
            in3 => \N__19193\,
            lcout => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19688\,
            in2 => \_gnd_net_\,
            in3 => \N__19190\,
            lcout => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__20867\,
            in1 => \N__19856\,
            in2 => \N__20714\,
            in3 => \N__19187\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__21035\,
            in1 => \N__21054\,
            in2 => \N__20600\,
            in3 => \N__20702\,
            lcout => \pwm_generator_inst.un19_threshold_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__20703\,
            in1 => \N__21020\,
            in2 => \N__20123\,
            in3 => \N__20996\,
            lcout => \pwm_generator_inst.un19_threshold_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_axb_4_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19427\,
            in2 => \N__19409\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19394\,
            in2 => \N__19376\,
            in3 => \N__19361\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19358\,
            in2 => \N__19343\,
            in3 => \N__19328\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19325\,
            in2 => \N__19307\,
            in3 => \N__19292\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19289\,
            in2 => \N__19271\,
            in3 => \N__19253\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19250\,
            in2 => \N__19232\,
            in3 => \N__19214\,
            lcout => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19670\,
            in2 => \N__19652\,
            in3 => \N__19637\,
            lcout => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19634\,
            in2 => \N__19616\,
            in3 => \N__19601\,
            lcout => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19598\,
            in2 => \N__19580\,
            in3 => \N__19565\,
            lcout => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \bfn_1_20_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19562\,
            in2 => \N__19544\,
            in3 => \N__19529\,
            lcout => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19526\,
            in2 => \N__19807\,
            in3 => \N__19511\,
            lcout => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19793\,
            in2 => \N__19508\,
            in3 => \N__19487\,
            lcout => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19484\,
            in2 => \N__19808\,
            in3 => \N__19466\,
            lcout => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19797\,
            in2 => \N__19463\,
            in3 => \N__19442\,
            lcout => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19844\,
            in2 => \N__19809\,
            in3 => \N__19826\,
            lcout => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19801\,
            in2 => \N__19763\,
            in3 => \N__19748\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19745\,
            in1 => \N__20054\,
            in2 => \_gnd_net_\,
            in3 => \N__19736\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\,
            ltout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__20723\,
            in1 => \N__20194\,
            in2 => \N__19733\,
            in3 => \N__20747\,
            lcout => \pwm_generator_inst.un19_threshold_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__20981\,
            in1 => \N__20954\,
            in2 => \N__20708\,
            in3 => \N__20504\,
            lcout => \pwm_generator_inst.un19_threshold_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20578\,
            in1 => \N__20921\,
            in2 => \N__20945\,
            in3 => \N__20695\,
            lcout => \pwm_generator_inst.un19_threshold_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__20912\,
            in1 => \N__21164\,
            in2 => \N__20709\,
            in3 => \N__21176\,
            lcout => \pwm_generator_inst.un19_threshold_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__20690\,
            in1 => \N__21128\,
            in2 => \N__21146\,
            in3 => \N__20882\,
            lcout => \pwm_generator_inst.un19_threshold_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011110000100"
        )
    port map (
            in0 => \N__21086\,
            in1 => \N__20689\,
            in2 => \N__20900\,
            in3 => \N__21098\,
            lcout => \pwm_generator_inst.un19_threshold_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20632\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_22_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19961\,
            in2 => \_gnd_net_\,
            in3 => \N__19952\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19949\,
            in2 => \_gnd_net_\,
            in3 => \N__19940\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19937\,
            in2 => \_gnd_net_\,
            in3 => \N__19928\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19925\,
            in2 => \_gnd_net_\,
            in3 => \N__19913\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44716\,
            in2 => \N__19910\,
            in3 => \N__19898\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19895\,
            in2 => \N__44746\,
            in3 => \N__19886\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44720\,
            in2 => \N__19883\,
            in3 => \N__19871\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19868\,
            in2 => \_gnd_net_\,
            in3 => \N__20039\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\,
            ltout => OPEN,
            carryin => \bfn_1_23_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20036\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20024\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20015\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20006\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19997\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19988\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19979\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19970\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_24_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20084\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20075\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20066\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20057\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.N_86_i_i_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__30008\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49270\,
            lcout => \N_86_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__25508\,
            in1 => \N__23468\,
            in2 => \N__22316\,
            in3 => \N__23276\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50032\,
            ce => 'H',
            sr => \N__49211\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000001010001"
        )
    port map (
            in0 => \N__25509\,
            in1 => \N__23469\,
            in2 => \N__21938\,
            in3 => \N__23277\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50032\,
            ce => 'H',
            sr => \N__49211\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__25510\,
            in1 => \N__23467\,
            in2 => \N__22160\,
            in3 => \N__23269\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50021\,
            ce => 'H',
            sr => \N__49216\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21516\,
            in2 => \_gnd_net_\,
            in3 => \N__21234\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__21447\,
            in1 => \N__21489\,
            in2 => \N__20174\,
            in3 => \N__21195\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20096\,
            in1 => \N__21358\,
            in2 => \N__20171\,
            in3 => \N__21397\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24453\,
            in1 => \N__24725\,
            in2 => \N__24571\,
            in3 => \N__24678\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001111"
        )
    port map (
            in0 => \N__21592\,
            in1 => \N__20129\,
            in2 => \N__20563\,
            in3 => \N__20338\,
            lcout => \pwm_generator_inst.un14_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__21015\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20119\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001111"
        )
    port map (
            in0 => \N__21593\,
            in1 => \N__20102\,
            in2 => \N__20564\,
            in3 => \N__20339\,
            lcout => \pwm_generator_inst.un14_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21645\,
            in1 => \N__21276\,
            in2 => \_gnd_net_\,
            in3 => \N__21318\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__21590\,
            in1 => \N__20090\,
            in2 => \N__20562\,
            in3 => \N__20337\,
            lcout => \pwm_generator_inst.threshold_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__20336\,
            in1 => \N__21591\,
            in2 => \N__20414\,
            in3 => \N__20553\,
            lcout => \pwm_generator_inst.threshold_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__21589\,
            in1 => \N__20405\,
            in2 => \N__20561\,
            in3 => \N__20335\,
            lcout => \pwm_generator_inst.threshold_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__20529\,
            in1 => \N__20399\,
            in2 => \N__20364\,
            in3 => \N__21585\,
            lcout => \pwm_generator_inst.threshold_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__21587\,
            in1 => \N__20531\,
            in2 => \N__20393\,
            in3 => \N__20357\,
            lcout => \pwm_generator_inst.threshold_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__20532\,
            in1 => \N__21588\,
            in2 => \N__20366\,
            in3 => \N__20384\,
            lcout => \pwm_generator_inst.threshold_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__20530\,
            in1 => \N__20378\,
            in2 => \N__20365\,
            in3 => \N__21586\,
            lcout => \pwm_generator_inst.un14_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001111"
        )
    port map (
            in0 => \N__21584\,
            in1 => \N__20372\,
            in2 => \N__20560\,
            in3 => \N__20361\,
            lcout => \pwm_generator_inst.un14_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24564\,
            in2 => \_gnd_net_\,
            in3 => \N__24726\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__24104\,
            in1 => \N__23847\,
            in2 => \_gnd_net_\,
            in3 => \N__23931\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20198\,
            in2 => \_gnd_net_\,
            in3 => \N__20745\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20596\,
            in2 => \_gnd_net_\,
            in3 => \N__21055\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20943\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20579\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001101"
        )
    port map (
            in0 => \N__21744\,
            in1 => \N__21875\,
            in2 => \N__21797\,
            in3 => \N__21107\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20976\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20503\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20474\,
            in2 => \_gnd_net_\,
            in3 => \N__20486\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_2_21_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20456\,
            in2 => \_gnd_net_\,
            in3 => \N__20468\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20438\,
            in2 => \_gnd_net_\,
            in3 => \N__20450\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20432\,
            in1 => \N__20420\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20843\,
            in2 => \_gnd_net_\,
            in3 => \N__20855\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20825\,
            in2 => \_gnd_net_\,
            in3 => \N__20837\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20807\,
            in2 => \_gnd_net_\,
            in3 => \N__20819\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20789\,
            in2 => \_gnd_net_\,
            in3 => \N__20801\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20771\,
            in2 => \_gnd_net_\,
            in3 => \N__20783\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_2_22_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20753\,
            in2 => \_gnd_net_\,
            in3 => \N__20765\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20746\,
            in2 => \_gnd_net_\,
            in3 => \N__20717\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__20691\,
            in1 => \N__20636\,
            in2 => \_gnd_net_\,
            in3 => \N__20603\,
            lcout => \pwm_generator_inst.un19_threshold_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21059\,
            in3 => \N__21023\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21016\,
            in2 => \_gnd_net_\,
            in3 => \N__20984\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20977\,
            in2 => \_gnd_net_\,
            in3 => \N__20948\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20944\,
            in2 => \_gnd_net_\,
            in3 => \N__20915\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21159\,
            in2 => \_gnd_net_\,
            in3 => \N__20903\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_23_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21081\,
            in2 => \_gnd_net_\,
            in3 => \N__20885\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21120\,
            in2 => \_gnd_net_\,
            in3 => \N__20873\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20870\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21160\,
            in2 => \_gnd_net_\,
            in3 => \N__21175\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__21121\,
            in1 => \_gnd_net_\,
            in2 => \N__21145\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__22588\,
            in1 => \N__22558\,
            in2 => \_gnd_net_\,
            in3 => \N__26027\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21082\,
            in2 => \_gnd_net_\,
            in3 => \N__21097\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.un7_start_stop_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__30007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49269\,
            lcout => un7_start_stop,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100000001"
        )
    port map (
            in0 => \N__23270\,
            in1 => \N__25479\,
            in2 => \N__23474\,
            in3 => \N__22232\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50033\,
            ce => 'H',
            sr => \N__49204\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__21989\,
            in1 => \N__23453\,
            in2 => \_gnd_net_\,
            in3 => \N__23272\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50033\,
            ce => 'H',
            sr => \N__49204\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001011001000"
        )
    port map (
            in0 => \N__23271\,
            in1 => \N__22039\,
            in2 => \N__23475\,
            in3 => \N__23660\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50033\,
            ce => 'H',
            sr => \N__49204\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101010"
        )
    port map (
            in0 => \N__25512\,
            in1 => \N__22094\,
            in2 => \N__23476\,
            in3 => \N__23274\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50022\,
            ce => 'H',
            sr => \N__49208\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000010110001"
        )
    port map (
            in0 => \N__23273\,
            in1 => \N__25514\,
            in2 => \N__22208\,
            in3 => \N__23466\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50022\,
            ce => 'H',
            sr => \N__49208\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001000101"
        )
    port map (
            in0 => \N__25513\,
            in1 => \N__21887\,
            in2 => \N__23477\,
            in3 => \N__23275\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50022\,
            ce => 'H',
            sr => \N__49208\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001111100000"
        )
    port map (
            in0 => \N__23436\,
            in1 => \N__23264\,
            in2 => \N__22073\,
            in3 => \N__25522\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50011\,
            ce => 'H',
            sr => \N__49212\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__25521\,
            in1 => \N__23437\,
            in2 => \N__23285\,
            in3 => \N__22298\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50011\,
            ce => 'H',
            sr => \N__49212\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011011000"
        )
    port map (
            in0 => \N__23258\,
            in1 => \N__21968\,
            in2 => \N__25523\,
            in3 => \N__23423\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50000\,
            ce => 'H',
            sr => \N__49217\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23420\,
            in1 => \N__25516\,
            in2 => \N__22289\,
            in3 => \N__23262\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50000\,
            ce => 'H',
            sr => \N__49217\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__25515\,
            in1 => \N__23422\,
            in2 => \N__23284\,
            in3 => \N__22271\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50000\,
            ce => 'H',
            sr => \N__49217\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23421\,
            in1 => \N__25517\,
            in2 => \N__22262\,
            in3 => \N__23263\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50000\,
            ce => 'H',
            sr => \N__49217\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21218\,
            in2 => \N__21254\,
            in3 => \N__21242\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_3_16_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21545\,
            in2 => \N__21212\,
            in3 => \N__21200\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21500\,
            in2 => \N__21536\,
            in3 => \N__21524\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21494\,
            in1 => \N__21458\,
            in2 => \N__21470\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21452\,
            in1 => \N__21419\,
            in2 => \N__21428\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21377\,
            in2 => \N__21413\,
            in3 => \N__21401\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21338\,
            in2 => \N__21371\,
            in3 => \N__21362\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21299\,
            in2 => \N__21332\,
            in3 => \N__21323\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21260\,
            in2 => \N__21293\,
            in3 => \N__21284\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_3_17_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21629\,
            in2 => \N__21662\,
            in3 => \N__21653\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21623\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49979\,
            ce => 'H',
            sr => \N__49228\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23848\,
            in1 => \N__23932\,
            in2 => \N__24028\,
            in3 => \N__23796\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__24115\,
            in1 => \N__24197\,
            in2 => \N__21596\,
            in3 => \N__24276\,
            lcout => \current_shift_inst.PI_CTRL.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30421\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49964\,
            ce => 'H',
            sr => \N__49237\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30199\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49964\,
            ce => 'H',
            sr => \N__49237\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30133\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49964\,
            ce => 'H',
            sr => \N__49237\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30481\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49964\,
            ce => 'H',
            sr => \N__49237\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__21793\,
            in1 => \N__21745\,
            in2 => \N__21719\,
            in3 => \N__21866\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22508\,
            in1 => \N__22625\,
            in2 => \N__22502\,
            in3 => \N__22514\,
            lcout => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\,
            ltout => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25235\,
            in2 => \N__21689\,
            in3 => \N__21674\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23973\,
            in2 => \_gnd_net_\,
            in3 => \N__25180\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25179\,
            in2 => \_gnd_net_\,
            in3 => \N__24066\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__23974\,
            in1 => \N__25353\,
            in2 => \N__21686\,
            in3 => \N__23901\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => \current_shift_inst.PI_CTRL.N_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__25236\,
            in1 => \N__24157\,
            in2 => \N__21683\,
            in3 => \N__25269\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23902\,
            in1 => \N__21680\,
            in2 => \N__24071\,
            in3 => \N__25354\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__25268\,
            in1 => \N__24156\,
            in2 => \N__25240\,
            in3 => \N__21673\,
            lcout => \current_shift_inst.PI_CTRL.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22056\,
            in2 => \_gnd_net_\,
            in3 => \N__21708\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__25317\,
            in1 => \N__21837\,
            in2 => \N__21878\,
            in3 => \N__25108\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25109\,
            in1 => \N__25318\,
            in2 => \N__21844\,
            in3 => \N__22057\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24155\,
            in2 => \_gnd_net_\,
            in3 => \N__24237\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__21808\,
            in1 => \N__25227\,
            in2 => \N__21857\,
            in3 => \N__25139\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => \current_shift_inst.PI_CTRL.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__21763\,
            in1 => \N__21854\,
            in2 => \N__21848\,
            in3 => \N__24238\,
            lcout => \current_shift_inst.PI_CTRL.N_160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000100"
        )
    port map (
            in0 => \N__25241\,
            in1 => \N__23975\,
            in2 => \N__25152\,
            in3 => \N__25281\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49246\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__24158\,
            in1 => \N__21821\,
            in2 => \N__21812\,
            in3 => \N__25147\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49246\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__24239\,
            in1 => \N__21764\,
            in2 => \_gnd_net_\,
            in3 => \N__21752\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49246\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100100010"
        )
    port map (
            in0 => \N__25280\,
            in1 => \N__25243\,
            in2 => \N__25154\,
            in3 => \N__24070\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49246\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000100"
        )
    port map (
            in0 => \N__25242\,
            in1 => \N__23903\,
            in2 => \N__25153\,
            in3 => \N__25282\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49246\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29126\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50046\,
            ce => 'H',
            sr => \N__49183\
        );

    \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23651\,
            in2 => \N__22040\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22019\,
            in2 => \N__23613\,
            in3 => \N__22007\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24255\,
            in2 => \N__22004\,
            in3 => \N__21983\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21980\,
            in2 => \N__24208\,
            in3 => \N__21956\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24111\,
            in2 => \N__21953\,
            in3 => \N__21923\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24003\,
            in2 => \N__21920\,
            in3 => \N__21905\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23921\,
            in2 => \N__21902\,
            in3 => \N__21881\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23834\,
            in2 => \N__22250\,
            in3 => \N__22226\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23789\,
            in2 => \N__22223\,
            in3 => \N__22199\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23736\,
            in2 => \N__22196\,
            in3 => \N__22181\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24733\,
            in2 => \N__22178\,
            in3 => \N__22145\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22142\,
            in2 => \N__24668\,
            in3 => \N__22130\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24614\,
            in2 => \N__22127\,
            in3 => \N__22112\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24551\,
            in2 => \N__22109\,
            in3 => \N__22088\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22085\,
            in2 => \N__24500\,
            in3 => \N__22064\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24446\,
            in2 => \N__22784\,
            in3 => \N__22304\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24396\,
            in2 => \N__22733\,
            in3 => \N__22301\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24329\,
            in2 => \N__22682\,
            in3 => \N__22292\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22637\,
            in2 => \N__25065\,
            in3 => \N__22280\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25010\,
            in2 => \N__23093\,
            in3 => \N__22277\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24962\,
            in2 => \N__23057\,
            in3 => \N__22274\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24911\,
            in2 => \N__23021\,
            in3 => \N__22265\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22988\,
            in2 => \N__24865\,
            in3 => \N__22253\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24814\,
            in2 => \N__22955\,
            in3 => \N__22352\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25877\,
            in2 => \N__22922\,
            in3 => \N__22349\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_4_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22886\,
            in2 => \N__25996\,
            in3 => \N__22346\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25953\,
            in2 => \N__22862\,
            in3 => \N__22343\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25914\,
            in2 => \N__23576\,
            in3 => \N__22340\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25617\,
            in2 => \N__23540\,
            in3 => \N__22337\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25563\,
            in2 => \N__23507\,
            in3 => \N__22334\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27032\,
            in1 => \N__25408\,
            in2 => \N__23492\,
            in3 => \N__22331\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23425\,
            in1 => \N__25505\,
            in2 => \N__22328\,
            in3 => \N__23181\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => 'H',
            sr => \N__49218\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__25503\,
            in1 => \N__23429\,
            in2 => \N__23222\,
            in3 => \N__22439\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => 'H',
            sr => \N__49218\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23424\,
            in1 => \N__25507\,
            in2 => \N__22433\,
            in3 => \N__23168\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => 'H',
            sr => \N__49218\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__25501\,
            in1 => \N__23427\,
            in2 => \N__23220\,
            in3 => \N__22421\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => 'H',
            sr => \N__49218\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23426\,
            in1 => \N__25506\,
            in2 => \N__22415\,
            in3 => \N__23182\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => 'H',
            sr => \N__49218\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__25504\,
            in1 => \N__23430\,
            in2 => \N__23223\,
            in3 => \N__22406\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => 'H',
            sr => \N__49218\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__25502\,
            in1 => \N__23428\,
            in2 => \N__23221\,
            in3 => \N__22400\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => 'H',
            sr => \N__49218\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22379\,
            in1 => \N__22358\,
            in2 => \N__22394\,
            in3 => \N__22478\,
            lcout => \current_shift_inst.PI_CTRL.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25616\,
            in1 => \N__24628\,
            in2 => \N__24508\,
            in3 => \N__23757\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__23806\,
            in1 => \N__22472\,
            in2 => \N__22373\,
            in3 => \N__24029\,
            lcout => \current_shift_inst.PI_CTRL.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25064\,
            in1 => \N__24916\,
            in2 => \N__24400\,
            in3 => \N__24333\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__25404\,
            in1 => \N__24864\,
            in2 => \N__22481\,
            in3 => \N__23702\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000111"
        )
    port map (
            in0 => \N__24277\,
            in1 => \N__23623\,
            in2 => \N__24207\,
            in3 => \N__23673\,
            lcout => \current_shift_inst.PI_CTRL.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24501\,
            in1 => \N__24627\,
            in2 => \N__23761\,
            in3 => \N__24454\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24679\,
            in1 => \N__22466\,
            in2 => \N__22457\,
            in3 => \N__25567\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24915\,
            in1 => \N__24337\,
            in2 => \N__25069\,
            in3 => \N__24392\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25618\,
            in1 => \N__24863\,
            in2 => \N__22454\,
            in3 => \N__22451\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23690\,
            in2 => \_gnd_net_\,
            in3 => \N__23674\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49955\,
            ce => 'H',
            sr => \N__49234\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23723\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24640\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25643\,
            in1 => \N__24695\,
            in2 => \N__22442\,
            in3 => \N__22619\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24418\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24469\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23722\,
            in1 => \N__25592\,
            in2 => \N__24419\,
            in3 => \N__24470\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24641\,
            in1 => \N__24694\,
            in2 => \N__22517\,
            in3 => \N__22493\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24833\,
            in1 => \N__24787\,
            in2 => \N__24593\,
            in3 => \N__24526\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24772\,
            in1 => \N__24985\,
            in2 => \N__24757\,
            in3 => \N__25030\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25031\,
            in1 => \N__24527\,
            in2 => \N__24989\,
            in3 => \N__24592\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24304\,
            in2 => \_gnd_net_\,
            in3 => \N__24358\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24887\,
            in1 => \N__24773\,
            in2 => \N__24761\,
            in3 => \N__22487\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24886\,
            in2 => \_gnd_net_\,
            in3 => \N__24937\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25661\,
            in1 => \N__25639\,
            in2 => \N__22628\,
            in3 => \N__25537\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25588\,
            in1 => \N__24832\,
            in2 => \N__24788\,
            in3 => \N__24938\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25660\,
            in1 => \N__24305\,
            in2 => \N__24362\,
            in3 => \N__25538\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22613\,
            in1 => \N__22604\,
            in2 => \N__22598\,
            in3 => \N__22595\,
            lcout => \current_shift_inst.PI_CTRL.N_158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25082\,
            in2 => \_gnd_net_\,
            in3 => \N__26040\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49244\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26041\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22568\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49244\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__22538\,
            in1 => \N__23438\,
            in2 => \_gnd_net_\,
            in3 => \N__23268\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50012\,
            ce => 'H',
            sr => \N__49194\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__23281\,
            in1 => \N__25475\,
            in2 => \N__23473\,
            in3 => \N__22532\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49200\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000001010001"
        )
    port map (
            in0 => \N__25471\,
            in1 => \N__23440\,
            in2 => \N__22526\,
            in3 => \N__23283\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49200\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__23278\,
            in1 => \N__25472\,
            in2 => \N__23470\,
            in3 => \N__22850\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49200\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__23280\,
            in1 => \N__25474\,
            in2 => \N__23472\,
            in3 => \N__22844\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49200\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__25470\,
            in1 => \N__23439\,
            in2 => \N__22838\,
            in3 => \N__23282\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49200\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__23279\,
            in1 => \N__25473\,
            in2 => \N__23471\,
            in3 => \N__22829\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49200\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22823\,
            in2 => \N__22808\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_16\,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22772\,
            in2 => \N__22751\,
            in3 => \N__22724\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22721\,
            in2 => \N__22700\,
            in3 => \N__22673\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22670\,
            in2 => \N__22652\,
            in3 => \N__22631\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23108\,
            in2 => \N__27110\,
            in3 => \N__23081\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23078\,
            in2 => \N__27112\,
            in3 => \N__23045\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23042\,
            in2 => \N__27111\,
            in3 => \N__23012\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23009\,
            in2 => \N__27113\,
            in3 => \N__22982\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27090\,
            in2 => \N__22979\,
            in3 => \N__22946\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_24\,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22943\,
            in2 => \N__27114\,
            in3 => \N__22913\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27094\,
            in2 => \N__22910\,
            in3 => \N__22880\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22877\,
            in2 => \N__27115\,
            in3 => \N__22853\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23591\,
            in2 => \N__27120\,
            in3 => \N__23564\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23561\,
            in2 => \N__27116\,
            in3 => \N__23531\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23528\,
            in2 => \N__27121\,
            in3 => \N__23498\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23495\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23385\,
            in1 => \N__25435\,
            in2 => \N__23224\,
            in3 => \N__23483\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49970\,
            ce => 'H',
            sr => \N__49213\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23386\,
            in1 => \N__25436\,
            in2 => \N__23225\,
            in3 => \N__23309\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49970\,
            ce => 'H',
            sr => \N__49213\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23696\,
            in1 => \N__23303\,
            in2 => \N__25850\,
            in3 => \N__23291\,
            lcout => \current_shift_inst.PI_CTRL.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25910\,
            in1 => \N__25949\,
            in2 => \N__25881\,
            in3 => \N__25559\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25985\,
            in2 => \_gnd_net_\,
            in3 => \N__24963\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24806\,
            in1 => \N__25011\,
            in2 => \N__23711\,
            in3 => \N__23708\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25012\,
            in1 => \N__24807\,
            in2 => \N__24974\,
            in3 => \N__25403\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30166\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49956\,
            ce => 'H',
            sr => \N__49223\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30106\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49956\,
            ce => 'H',
            sr => \N__49223\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30452\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49956\,
            ce => 'H',
            sr => \N__49223\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30070\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49956\,
            ce => 'H',
            sr => \N__49223\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23689\,
            in2 => \N__23675\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23630\,
            in2 => \N__23624\,
            in3 => \N__23594\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49229\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24290\,
            in2 => \N__24281\,
            in3 => \N__24218\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49229\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24215\,
            in2 => \N__24209\,
            in3 => \N__24125\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49229\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24122\,
            in2 => \N__24116\,
            in3 => \N__24032\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49229\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24024\,
            in2 => \N__23987\,
            in3 => \N__23948\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49229\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23945\,
            in2 => \N__23939\,
            in3 => \N__23867\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49229\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23864\,
            in2 => \N__23855\,
            in3 => \N__23813\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49229\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25802\,
            in2 => \N__23810\,
            in3 => \N__23765\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_5_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__49941\,
            ce => 'H',
            sr => \N__49235\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26273\,
            in2 => \N__23762\,
            in3 => \N__23714\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__49941\,
            ce => 'H',
            sr => \N__49235\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25823\,
            in2 => \N__24740\,
            in3 => \N__24686\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__49941\,
            ce => 'H',
            sr => \N__49235\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26264\,
            in2 => \N__24683\,
            in3 => \N__24632\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__49941\,
            ce => 'H',
            sr => \N__49235\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25814\,
            in2 => \N__24629\,
            in3 => \N__24578\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__49941\,
            ce => 'H',
            sr => \N__49235\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26282\,
            in2 => \N__24575\,
            in3 => \N__24518\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__49941\,
            ce => 'H',
            sr => \N__49235\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27020\,
            in2 => \N__24515\,
            in3 => \N__24461\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__49941\,
            ce => 'H',
            sr => \N__49235\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24458\,
            in2 => \N__27839\,
            in3 => \N__24407\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__49941\,
            ce => 'H',
            sr => \N__49235\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26246\,
            in2 => \N__24404\,
            in3 => \N__24347\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_5_21_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49238\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26993\,
            in2 => \N__24344\,
            in3 => \N__24293\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49238\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26255\,
            in2 => \N__25076\,
            in3 => \N__25022\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49238\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27011\,
            in2 => \N__25019\,
            in3 => \N__24977\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49238\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27002\,
            in2 => \N__24973\,
            in3 => \N__24929\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49238\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27827\,
            in2 => \N__24926\,
            in3 => \N__24878\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49238\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26237\,
            in2 => \N__24875\,
            in3 => \N__24824\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49238\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29057\,
            in2 => \N__24821\,
            in3 => \N__24776\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49238\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27947\,
            in2 => \N__25889\,
            in3 => \N__24764\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_5_22_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49239\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27818\,
            in2 => \N__26000\,
            in3 => \N__25664\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49239\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26984\,
            in2 => \N__25964\,
            in3 => \N__25646\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49239\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29030\,
            in2 => \N__25928\,
            in3 => \N__25628\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49239\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29048\,
            in2 => \N__25625\,
            in3 => \N__25577\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49239\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29039\,
            in2 => \N__25574\,
            in3 => \N__25526\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49239\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27956\,
            in1 => \N__25511\,
            in2 => \_gnd_net_\,
            in3 => \N__25358\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49239\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__25214\,
            in1 => \N__25140\,
            in2 => \N__25355\,
            in3 => \N__25288\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49923\,
            ce => 'H',
            sr => \N__49240\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__25289\,
            in1 => \N__25215\,
            in2 => \N__25181\,
            in3 => \N__25151\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49923\,
            ce => 'H',
            sr => \N__49240\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25835\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49923\,
            ce => 'H',
            sr => \N__49240\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__28820\,
            in1 => \N__25708\,
            in2 => \_gnd_net_\,
            in3 => \N__29118\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => \phase_controller_inst2.stoper_tr.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101011111010"
        )
    port map (
            in0 => \N__25709\,
            in1 => \N__28747\,
            in2 => \N__25712\,
            in3 => \N__28821\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50023\,
            ce => 'H',
            sr => \N__49168\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28766\,
            in2 => \_gnd_net_\,
            in3 => \N__26221\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28819\,
            in2 => \_gnd_net_\,
            in3 => \N__28743\,
            lcout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25700\,
            in3 => \N__28767\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26456\,
            in2 => \N__25697\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26196\,
            in1 => \N__26414\,
            in2 => \_gnd_net_\,
            in3 => \N__25685\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__50013\,
            ce => 'H',
            sr => \N__49173\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__26204\,
            in1 => \N__26381\,
            in2 => \N__25682\,
            in3 => \N__25670\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__50013\,
            ce => 'H',
            sr => \N__49173\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26197\,
            in1 => \N__26348\,
            in2 => \_gnd_net_\,
            in3 => \N__25667\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__50013\,
            ce => 'H',
            sr => \N__49173\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26205\,
            in1 => \N__26672\,
            in2 => \_gnd_net_\,
            in3 => \N__25739\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__50013\,
            ce => 'H',
            sr => \N__49173\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26198\,
            in1 => \N__26651\,
            in2 => \_gnd_net_\,
            in3 => \N__25736\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__50013\,
            ce => 'H',
            sr => \N__49173\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26206\,
            in1 => \N__26618\,
            in2 => \_gnd_net_\,
            in3 => \N__25733\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__50013\,
            ce => 'H',
            sr => \N__49173\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26199\,
            in1 => \N__26597\,
            in2 => \_gnd_net_\,
            in3 => \N__25730\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__50013\,
            ce => 'H',
            sr => \N__49173\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26203\,
            in1 => \N__26570\,
            in2 => \_gnd_net_\,
            in3 => \N__25727\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__50002\,
            ce => 'H',
            sr => \N__49179\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26192\,
            in1 => \N__26537\,
            in2 => \_gnd_net_\,
            in3 => \N__25724\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__50002\,
            ce => 'H',
            sr => \N__49179\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26200\,
            in1 => \N__26519\,
            in2 => \_gnd_net_\,
            in3 => \N__25721\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__50002\,
            ce => 'H',
            sr => \N__49179\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26193\,
            in1 => \N__26489\,
            in2 => \_gnd_net_\,
            in3 => \N__25718\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__50002\,
            ce => 'H',
            sr => \N__49179\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26201\,
            in1 => \N__26768\,
            in2 => \_gnd_net_\,
            in3 => \N__25715\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__50002\,
            ce => 'H',
            sr => \N__49179\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26194\,
            in1 => \N__26749\,
            in2 => \_gnd_net_\,
            in3 => \N__25766\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__50002\,
            ce => 'H',
            sr => \N__49179\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26202\,
            in1 => \N__26723\,
            in2 => \_gnd_net_\,
            in3 => \N__25763\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__50002\,
            ce => 'H',
            sr => \N__49179\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26195\,
            in1 => \N__27211\,
            in2 => \_gnd_net_\,
            in3 => \N__25760\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__50002\,
            ce => 'H',
            sr => \N__49179\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26173\,
            in1 => \N__27238\,
            in2 => \_gnd_net_\,
            in3 => \N__25757\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__49989\,
            ce => 'H',
            sr => \N__49184\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26177\,
            in1 => \N__26298\,
            in2 => \_gnd_net_\,
            in3 => \N__25754\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__49989\,
            ce => 'H',
            sr => \N__49184\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26174\,
            in1 => \N__26319\,
            in2 => \_gnd_net_\,
            in3 => \N__25751\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__49989\,
            ce => 'H',
            sr => \N__49184\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26178\,
            in1 => \N__26842\,
            in2 => \_gnd_net_\,
            in3 => \N__25748\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__49989\,
            ce => 'H',
            sr => \N__49184\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26175\,
            in1 => \N__26824\,
            in2 => \_gnd_net_\,
            in3 => \N__25745\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__49989\,
            ce => 'H',
            sr => \N__49184\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26179\,
            in1 => \N__27321\,
            in2 => \_gnd_net_\,
            in3 => \N__25742\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__49989\,
            ce => 'H',
            sr => \N__49184\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26176\,
            in1 => \N__27295\,
            in2 => \_gnd_net_\,
            in3 => \N__25793\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__49989\,
            ce => 'H',
            sr => \N__49184\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26180\,
            in1 => \N__27744\,
            in2 => \_gnd_net_\,
            in3 => \N__25790\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__49989\,
            ce => 'H',
            sr => \N__49184\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26169\,
            in1 => \N__27777\,
            in2 => \_gnd_net_\,
            in3 => \N__25787\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__49981\,
            ce => 'H',
            sr => \N__49189\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26207\,
            in1 => \N__26930\,
            in2 => \_gnd_net_\,
            in3 => \N__25784\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__49981\,
            ce => 'H',
            sr => \N__49189\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26170\,
            in1 => \N__26947\,
            in2 => \_gnd_net_\,
            in3 => \N__25781\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__49981\,
            ce => 'H',
            sr => \N__49189\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26208\,
            in1 => \N__27565\,
            in2 => \_gnd_net_\,
            in3 => \N__25778\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__49981\,
            ce => 'H',
            sr => \N__49189\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26171\,
            in1 => \N__27594\,
            in2 => \_gnd_net_\,
            in3 => \N__25775\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__49981\,
            ce => 'H',
            sr => \N__49189\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26209\,
            in1 => \N__27489\,
            in2 => \_gnd_net_\,
            in3 => \N__25772\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__49981\,
            ce => 'H',
            sr => \N__49189\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26172\,
            in1 => \N__27519\,
            in2 => \_gnd_net_\,
            in3 => \N__25769\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49981\,
            ce => 'H',
            sr => \N__49189\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__31235\,
            in1 => \N__31196\,
            in2 => \N__31167\,
            in3 => \N__32688\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49971\,
            ce => 'H',
            sr => \N__49195\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31954\,
            in2 => \_gnd_net_\,
            in3 => \N__38392\,
            lcout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26003\,
            in3 => \N__36696\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28834\,
            in2 => \_gnd_net_\,
            in3 => \N__29119\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25995\,
            in1 => \N__25957\,
            in2 => \N__25924\,
            in3 => \N__25882\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29632\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49936\,
            ce => 'H',
            sr => \N__49219\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30322\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49224\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30268\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49224\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30379\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49224\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30235\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49224\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30352\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49224\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30298\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49224\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30592\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49230\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30655\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49230\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30967\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49230\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36700\,
            in2 => \_gnd_net_\,
            in3 => \N__36724\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__28783\,
            in1 => \N__26228\,
            in2 => \N__26443\,
            in3 => \N__26181\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49916\,
            ce => 'H',
            sr => \N__49236\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26057\,
            in2 => \_gnd_net_\,
            in3 => \N__26045\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49916\,
            ce => 'H',
            sr => \N__49236\
        );

    \phase_controller_inst2.stoper_tr.target_time_28_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35370\,
            in1 => \N__28393\,
            in2 => \_gnd_net_\,
            in3 => \N__32411\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50040\,
            ce => \N__28913\,
            sr => \N__49146\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32357\,
            in1 => \N__29180\,
            in2 => \_gnd_net_\,
            in3 => \N__33838\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50034\,
            ce => \N__28914\,
            sr => \N__49153\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27188\,
            in1 => \N__34469\,
            in2 => \_gnd_net_\,
            in3 => \N__32330\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50024\,
            ce => \N__28915\,
            sr => \N__49158\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__32328\,
            in1 => \N__28044\,
            in2 => \N__34400\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50024\,
            ce => \N__28915\,
            sr => \N__49158\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28506\,
            in1 => \N__33617\,
            in2 => \_gnd_net_\,
            in3 => \N__32332\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50024\,
            ce => \N__28915\,
            sr => \N__49158\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33476\,
            in1 => \N__27173\,
            in2 => \_gnd_net_\,
            in3 => \N__32333\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50024\,
            ce => \N__28915\,
            sr => \N__49158\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32329\,
            in1 => \N__27270\,
            in2 => \_gnd_net_\,
            in3 => \N__35015\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50024\,
            ce => \N__28915\,
            sr => \N__49158\
        );

    \phase_controller_inst2.stoper_tr.target_time_23_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29417\,
            in1 => \N__34646\,
            in2 => \_gnd_net_\,
            in3 => \N__32331\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50024\,
            ce => \N__28915\,
            sr => \N__49158\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__26321\,
            in1 => \N__26299\,
            in2 => \N__26468\,
            in3 => \N__26330\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__26329\,
            in1 => \N__26320\,
            in2 => \N__26303\,
            in3 => \N__26464\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31076\,
            in1 => \N__34942\,
            in2 => \_gnd_net_\,
            in3 => \N__32405\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50014\,
            ce => \N__28916\,
            sr => \N__49163\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32404\,
            in1 => \N__29204\,
            in2 => \_gnd_net_\,
            in3 => \N__29240\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50014\,
            ce => \N__28916\,
            sr => \N__49163\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27988\,
            in1 => \N__33908\,
            in2 => \_gnd_net_\,
            in3 => \N__32406\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50014\,
            ce => \N__28916\,
            sr => \N__49163\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33768\,
            in1 => \N__28589\,
            in2 => \_gnd_net_\,
            in3 => \N__32407\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50014\,
            ce => \N__28916\,
            sr => \N__49163\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27374\,
            in2 => \N__26423\,
            in3 => \N__26455\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26413\,
            in1 => \N__26402\,
            in2 => \N__26396\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26387\,
            in2 => \N__26369\,
            in3 => \N__26380\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26336\,
            in2 => \N__26360\,
            in3 => \N__26347\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26678\,
            in2 => \N__26660\,
            in3 => \N__26671\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26777\,
            in2 => \N__26639\,
            in3 => \N__26650\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26627\,
            in2 => \N__26606\,
            in3 => \N__26617\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26585\,
            in2 => \N__26972\,
            in3 => \N__26596\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26579\,
            in2 => \N__26558\,
            in3 => \N__26569\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26525\,
            in2 => \N__26549\,
            in3 => \N__26536\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26518\,
            in1 => \N__26507\,
            in2 => \N__26498\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27644\,
            in2 => \N__26477\,
            in3 => \N__26488\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26756\,
            in2 => \N__27431\,
            in3 => \N__26767\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27422\,
            in2 => \N__26735\,
            in3 => \N__26750\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26711\,
            in2 => \N__27404\,
            in3 => \N__26722\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27251\,
            in2 => \N__27197\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26705\,
            in2 => \N__26693\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26852\,
            in2 => \N__26807\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27281\,
            in2 => \N__27368\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27158\,
            in2 => \N__27722\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26915\,
            in2 => \N__26960\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27530\,
            in2 => \N__26885\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27470\,
            in2 => \N__26870\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26855\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__26786\,
            in1 => \N__26795\,
            in2 => \N__26843\,
            in3 => \N__26823\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__26794\,
            in1 => \N__26841\,
            in2 => \N__26825\,
            in3 => \N__26785\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_20_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32359\,
            in1 => \N__27889\,
            in2 => \_gnd_net_\,
            in3 => \N__34852\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49972\,
            ce => \N__28919\,
            sr => \N__49185\
        );

    \phase_controller_inst2.stoper_tr.target_time_21_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34784\,
            in1 => \N__31310\,
            in2 => \_gnd_net_\,
            in3 => \N__32362\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49972\,
            ce => \N__28919\,
            sr => \N__49185\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32360\,
            in1 => \N__28638\,
            in2 => \_gnd_net_\,
            in3 => \N__33689\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49972\,
            ce => \N__28919\,
            sr => \N__49185\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33544\,
            in1 => \N__28471\,
            in2 => \_gnd_net_\,
            in3 => \N__32358\,
            lcout => \elapsed_time_ns_1_RNIKJ91B_0_8\,
            ltout => \elapsed_time_ns_1_RNIKJ91B_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32361\,
            in1 => \_gnd_net_\,
            in2 => \N__26975\,
            in3 => \N__33545\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49972\,
            ce => \N__28919\,
            sr => \N__49185\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__26929\,
            in1 => \N__26906\,
            in2 => \N__26897\,
            in3 => \N__26946\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__26905\,
            in1 => \N__26896\,
            in2 => \N__26948\,
            in3 => \N__26928\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_26_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27860\,
            in1 => \N__35531\,
            in2 => \_gnd_net_\,
            in3 => \N__32421\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49965\,
            ce => \N__28921\,
            sr => \N__49190\
        );

    \phase_controller_inst2.stoper_tr.target_time_27_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32419\,
            in1 => \N__35441\,
            in2 => \_gnd_net_\,
            in3 => \N__27464\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49965\,
            ce => \N__28921\,
            sr => \N__49190\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__27623\,
            in1 => \N__27564\,
            in2 => \N__27598\,
            in3 => \N__27544\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_29_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32420\,
            in1 => \N__35276\,
            in2 => \_gnd_net_\,
            in3 => \N__28427\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49965\,
            ce => \N__28921\,
            sr => \N__49190\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011101111"
        )
    port map (
            in0 => \N__27679\,
            in1 => \N__27520\,
            in2 => \N__27496\,
            in3 => \N__27694\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__27709\,
            in1 => \N__27784\,
            in2 => \N__27757\,
            in3 => \N__28937\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27146\,
            in2 => \_gnd_net_\,
            in3 => \N__27125\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30721\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49925\,
            ce => 'H',
            sr => \N__49220\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30565\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49225\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30535\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49225\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30622\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49225\
        );

    \current_shift_inst.PI_CTRL.prop_term_27_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30844\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49912\,
            ce => 'H',
            sr => \N__49231\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27275\,
            in1 => \N__35014\,
            in2 => \_gnd_net_\,
            in3 => \N__32410\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50041\,
            ce => \N__32737\,
            sr => \N__49135\
        );

    \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34718\,
            in1 => \N__28027\,
            in2 => \_gnd_net_\,
            in3 => \N__32409\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50035\,
            ce => \N__28912\,
            sr => \N__49139\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32353\,
            in1 => \N__34467\,
            in2 => \_gnd_net_\,
            in3 => \N__27187\,
            lcout => \elapsed_time_ns_1_RNIT6OBB_0_10\,
            ltout => \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__34468\,
            in1 => \_gnd_net_\,
            in2 => \N__27176\,
            in3 => \N__32355\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50025\,
            ce => \N__32738\,
            sr => \N__49147\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33474\,
            in1 => \N__27172\,
            in2 => \_gnd_net_\,
            in3 => \N__32352\,
            lcout => \elapsed_time_ns_1_RNILK91B_0_9\,
            ltout => \elapsed_time_ns_1_RNILK91B_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32354\,
            in1 => \_gnd_net_\,
            in2 => \N__27161\,
            in3 => \N__33475\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50025\,
            ce => \N__32738\,
            sr => \N__49147\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__27660\,
            in1 => \_gnd_net_\,
            in2 => \N__34319\,
            in3 => \N__32356\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50025\,
            ce => \N__32738\,
            sr => \N__49147\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32304\,
            in1 => \N__27664\,
            in2 => \_gnd_net_\,
            in3 => \N__34315\,
            lcout => \elapsed_time_ns_1_RNIV8OBB_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29271\,
            in1 => \N__27394\,
            in2 => \_gnd_net_\,
            in3 => \N__32307\,
            lcout => \elapsed_time_ns_1_RNIDC91B_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32306\,
            in1 => \N__28507\,
            in2 => \_gnd_net_\,
            in3 => \N__33616\,
            lcout => \elapsed_time_ns_1_RNIJI91B_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27989\,
            in1 => \N__33903\,
            in2 => \_gnd_net_\,
            in3 => \N__32308\,
            lcout => \elapsed_time_ns_1_RNIFE91B_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33902\,
            in1 => \N__29239\,
            in2 => \N__33839\,
            in3 => \N__29270\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31309\,
            in1 => \N__34776\,
            in2 => \_gnd_net_\,
            in3 => \N__32303\,
            lcout => \elapsed_time_ns_1_RNIV9PBB_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32309\,
            in1 => \N__28046\,
            in2 => \_gnd_net_\,
            in3 => \N__34396\,
            lcout => \elapsed_time_ns_1_RNIU7OBB_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27274\,
            in1 => \N__35007\,
            in2 => \_gnd_net_\,
            in3 => \N__32305\,
            lcout => \elapsed_time_ns_1_RNI5FOBB_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_20_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32397\,
            in1 => \_gnd_net_\,
            in2 => \N__27890\,
            in3 => \N__34856\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50003\,
            ce => \N__32721\,
            sr => \N__49159\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34101\,
            in1 => \N__27415\,
            in2 => \_gnd_net_\,
            in3 => \N__32394\,
            lcout => \elapsed_time_ns_1_RNI2COBB_0_15\,
            ltout => \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32395\,
            in1 => \_gnd_net_\,
            in2 => \N__27254\,
            in3 => \N__34102\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50003\,
            ce => \N__32721\,
            sr => \N__49159\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__27634\,
            in1 => \N__31871\,
            in2 => \N__31285\,
            in3 => \N__31901\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32396\,
            in1 => \N__27390\,
            in2 => \_gnd_net_\,
            in3 => \N__29272\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50003\,
            ce => \N__32721\,
            sr => \N__49159\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__27452\,
            in1 => \N__27220\,
            in2 => \N__27443\,
            in3 => \N__27245\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__27244\,
            in1 => \N__27451\,
            in2 => \N__27224\,
            in3 => \N__27439\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32400\,
            in1 => \N__29348\,
            in2 => \_gnd_net_\,
            in3 => \N__34044\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49990\,
            ce => \N__28917\,
            sr => \N__49164\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33974\,
            in1 => \N__32401\,
            in2 => \_gnd_net_\,
            in3 => \N__29381\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49990\,
            ce => \N__28917\,
            sr => \N__49164\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32398\,
            in1 => \_gnd_net_\,
            in2 => \N__29315\,
            in3 => \N__34244\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49990\,
            ce => \N__28917\,
            sr => \N__49164\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32006\,
            in1 => \N__34174\,
            in2 => \_gnd_net_\,
            in3 => \N__32402\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49990\,
            ce => \N__28917\,
            sr => \N__49164\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32399\,
            in1 => \N__34106\,
            in2 => \_gnd_net_\,
            in3 => \N__27416\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49990\,
            ce => \N__28917\,
            sr => \N__49164\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29273\,
            in1 => \N__27395\,
            in2 => \_gnd_net_\,
            in3 => \N__32403\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49990\,
            ce => \N__28917\,
            sr => \N__49164\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__27328\,
            in1 => \N__27347\,
            in2 => \N__27305\,
            in3 => \N__27359\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011101111"
        )
    port map (
            in0 => \N__27358\,
            in1 => \N__27346\,
            in2 => \N__27332\,
            in3 => \N__27304\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27668\,
            in1 => \N__34304\,
            in2 => \_gnd_net_\,
            in3 => \N__32408\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49982\,
            ce => \N__28918\,
            sr => \N__49169\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__27638\,
            in1 => \N__31870\,
            in2 => \N__31286\,
            in3 => \N__31900\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32393\,
            in1 => \N__33687\,
            in2 => \_gnd_net_\,
            in3 => \N__28639\,
            lcout => \elapsed_time_ns_1_RNIIH91B_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29307\,
            in1 => \N__32392\,
            in2 => \_gnd_net_\,
            in3 => \N__34239\,
            lcout => \elapsed_time_ns_1_RNI0AOBB_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__27622\,
            in1 => \N__27599\,
            in2 => \N__27572\,
            in3 => \N__27545\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__27524\,
            in1 => \N__27683\,
            in2 => \N__27500\,
            in3 => \N__27698\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011010100"
        )
    port map (
            in0 => \N__31712\,
            in1 => \N__27794\,
            in2 => \N__27806\,
            in3 => \N__31732\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__27793\,
            in1 => \N__31711\,
            in2 => \N__31736\,
            in3 => \N__27802\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35429\,
            in1 => \N__32417\,
            in2 => \_gnd_net_\,
            in3 => \N__27463\,
            lcout => \elapsed_time_ns_1_RNI5GPBB_0_27\,
            ltout => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_27_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__32418\,
            in1 => \N__35430\,
            in2 => \N__27809\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49966\,
            ce => \N__32679\,
            sr => \N__49180\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011101111"
        )
    port map (
            in0 => \N__32473\,
            in1 => \N__28666\,
            in2 => \N__32771\,
            in3 => \N__28654\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_26_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27859\,
            in1 => \N__35525\,
            in2 => \_gnd_net_\,
            in3 => \N__32426\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49957\,
            ce => \N__32560\,
            sr => \N__49186\
        );

    \phase_controller_inst1.stoper_tr.target_time_24_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32449\,
            in1 => \N__34577\,
            in2 => \_gnd_net_\,
            in3 => \N__32425\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49957\,
            ce => \N__32560\,
            sr => \N__49186\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__27710\,
            in1 => \N__27785\,
            in2 => \N__27758\,
            in3 => \N__28936\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_24_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__32453\,
            in1 => \N__32423\,
            in2 => \_gnd_net_\,
            in3 => \N__34576\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49948\,
            ce => \N__28922\,
            sr => \N__49191\
        );

    \phase_controller_inst2.stoper_tr.target_time_31_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35149\,
            in1 => \N__32424\,
            in2 => \_gnd_net_\,
            in3 => \N__28975\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49948\,
            ce => \N__28922\,
            sr => \N__49191\
        );

    \phase_controller_inst2.stoper_tr.target_time_30_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32422\,
            in1 => \N__28561\,
            in2 => \_gnd_net_\,
            in3 => \N__35192\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49948\,
            ce => \N__28922\,
            sr => \N__49191\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29807\,
            in2 => \_gnd_net_\,
            in3 => \N__31945\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27882\,
            in1 => \N__34845\,
            in2 => \_gnd_net_\,
            in3 => \N__32415\,
            lcout => \elapsed_time_ns_1_RNIU8PBB_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27858\,
            in1 => \N__35527\,
            in2 => \_gnd_net_\,
            in3 => \N__32416\,
            lcout => \elapsed_time_ns_1_RNI4FPBB_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101011001100"
        )
    port map (
            in0 => \N__31946\,
            in1 => \N__28866\,
            in2 => \N__38399\,
            in3 => \N__36692\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => 'H',
            sr => \N__49201\
        );

    \phase_controller_inst2.start_timer_hc_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__28847\,
            in1 => \N__28678\,
            in2 => \N__29813\,
            in3 => \N__33353\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => 'H',
            sr => \N__49201\
        );

    \phase_controller_inst2.state_2_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__29934\,
            in1 => \N__28883\,
            in2 => \N__29891\,
            in3 => \N__28867\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => 'H',
            sr => \N__49201\
        );

    \phase_controller_inst1.state_4_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__29995\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33352\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => 'H',
            sr => \N__49201\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29808\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => 'H',
            sr => \N__49201\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30691\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49214\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30508\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49221\
        );

    \current_shift_inst.PI_CTRL.prop_term_26_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30871\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49909\,
            ce => 'H',
            sr => \N__49226\
        );

    \current_shift_inst.PI_CTRL.prop_term_31_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30737\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49909\,
            ce => 'H',
            sr => \N__49226\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30901\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49909\,
            ce => 'H',
            sr => \N__49226\
        );

    \phase_controller_inst2.S1_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29887\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49895\,
            ce => 'H',
            sr => \N__49245\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27929\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31072\,
            in1 => \N__34943\,
            in2 => \_gnd_net_\,
            in3 => \N__32327\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50027\,
            ce => \N__32736\,
            sr => \N__49122\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__31534\,
            in1 => \N__27911\,
            in2 => \N__27902\,
            in3 => \N__31507\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__27910\,
            in1 => \N__31535\,
            in2 => \N__31508\,
            in3 => \N__27901\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32325\,
            in1 => \N__35374\,
            in2 => \_gnd_net_\,
            in3 => \N__28392\,
            lcout => \elapsed_time_ns_1_RNI6HPBB_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28028\,
            in1 => \N__34716\,
            in2 => \_gnd_net_\,
            in3 => \N__32326\,
            lcout => \elapsed_time_ns_1_RNI0BPBB_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_23_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34645\,
            in1 => \N__29412\,
            in2 => \_gnd_net_\,
            in3 => \N__32186\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__32702\,
            sr => \N__49136\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28045\,
            in1 => \N__34395\,
            in2 => \_gnd_net_\,
            in3 => \N__32185\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__32702\,
            sr => \N__49136\
        );

    \phase_controller_inst1.stoper_tr.target_time_22_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32184\,
            in1 => \N__28026\,
            in2 => \_gnd_net_\,
            in3 => \N__34717\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__32702\,
            sr => \N__49136\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29196\,
            in1 => \N__29229\,
            in2 => \_gnd_net_\,
            in3 => \N__32187\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__32702\,
            sr => \N__49136\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29175\,
            in1 => \N__33834\,
            in2 => \_gnd_net_\,
            in3 => \N__32188\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__32702\,
            sr => \N__49136\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__31843\,
            in1 => \N__28001\,
            in2 => \N__31819\,
            in3 => \N__28010\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__28009\,
            in1 => \N__28000\,
            in2 => \N__31820\,
            in3 => \N__31844\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27987\,
            in1 => \N__33907\,
            in2 => \_gnd_net_\,
            in3 => \N__32190\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49992\,
            ce => \N__32726\,
            sr => \N__49140\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27962\,
            in2 => \N__27971\,
            in3 => \N__31172\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28160\,
            in2 => \N__28151\,
            in3 => \N__31127\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28142\,
            in2 => \N__28136\,
            in3 => \N__31100\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28127\,
            in2 => \N__28118\,
            in3 => \N__31478\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28607\,
            in2 => \N__28109\,
            in3 => \N__31457\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31436\,
            in1 => \N__28100\,
            in2 => \N__28619\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28487\,
            in2 => \N__28094\,
            in3 => \N__31415\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28460\,
            in2 => \N__28085\,
            in3 => \N__31394\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28073\,
            in2 => \N__28064\,
            in3 => \N__31373\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28055\,
            in2 => \N__28283\,
            in3 => \N__31352\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28274\,
            in2 => \N__28262\,
            in3 => \N__31331\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28253\,
            in2 => \N__28241\,
            in3 => \N__31667\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29288\,
            in2 => \N__28232\,
            in3 => \N__31646\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28598\,
            in2 => \N__28223\,
            in3 => \N__31625\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28205\,
            in2 => \N__28214\,
            in3 => \N__31604\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29396\,
            in2 => \N__29390\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28199\,
            in2 => \N__28190\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28178\,
            in2 => \N__28172\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28352\,
            in2 => \N__28343\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28289\,
            in2 => \N__28520\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28328\,
            in2 => \N__28319\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28436\,
            in2 => \N__28448\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28361\,
            in2 => \N__28307\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28292\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__28544\,
            in1 => \N__31760\,
            in2 => \N__31787\,
            in3 => \N__28529\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_25_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28958\,
            in1 => \N__34508\,
            in2 => \_gnd_net_\,
            in3 => \N__32345\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49959\,
            ce => \N__32687\,
            sr => \N__49165\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__28543\,
            in1 => \N__31759\,
            in2 => \N__31786\,
            in3 => \N__28528\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32344\,
            in1 => \N__33609\,
            in2 => \_gnd_net_\,
            in3 => \N__28511\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49959\,
            ce => \N__32687\,
            sr => \N__49165\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33538\,
            in1 => \N__28478\,
            in2 => \_gnd_net_\,
            in3 => \N__32346\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49959\,
            ce => \N__32687\,
            sr => \N__49165\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__32792\,
            in1 => \N__31687\,
            in2 => \N__28406\,
            in3 => \N__28370\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__28369\,
            in1 => \N__32791\,
            in2 => \N__31691\,
            in3 => \N__28402\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35270\,
            in1 => \N__32338\,
            in2 => \_gnd_net_\,
            in3 => \N__28420\,
            lcout => \elapsed_time_ns_1_RNI7IPBB_0_29\,
            ltout => \elapsed_time_ns_1_RNI7IPBB_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_29_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32340\,
            in1 => \_gnd_net_\,
            in2 => \N__28409\,
            in3 => \N__35271\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49950\,
            ce => \N__32631\,
            sr => \N__49170\
        );

    \phase_controller_inst1.stoper_tr.target_time_28_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32339\,
            in1 => \N__35363\,
            in2 => \_gnd_net_\,
            in3 => \N__28394\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49950\,
            ce => \N__32631\,
            sr => \N__49170\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__32474\,
            in1 => \N__28667\,
            in2 => \N__32770\,
            in3 => \N__28655\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_30_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32347\,
            in1 => \N__28560\,
            in2 => \_gnd_net_\,
            in3 => \N__35191\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49943\,
            ce => \N__32627\,
            sr => \N__49174\
        );

    \phase_controller_inst1.stoper_tr.target_time_31_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32348\,
            in1 => \N__35148\,
            in2 => \_gnd_net_\,
            in3 => \N__28974\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49943\,
            ce => \N__32627\,
            sr => \N__49174\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33688\,
            in1 => \N__28643\,
            in2 => \_gnd_net_\,
            in3 => \N__32351\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49943\,
            ce => \N__32627\,
            sr => \N__49174\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32349\,
            in1 => \N__33770\,
            in2 => \_gnd_net_\,
            in3 => \N__28578\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49943\,
            ce => \N__32627\,
            sr => \N__49174\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32002\,
            in1 => \N__34175\,
            in2 => \_gnd_net_\,
            in3 => \N__32350\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49943\,
            ce => \N__32627\,
            sr => \N__49174\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32335\,
            in1 => \N__28957\,
            in2 => \_gnd_net_\,
            in3 => \N__34513\,
            lcout => \elapsed_time_ns_1_RNI3EPBB_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32334\,
            in1 => \N__33769\,
            in2 => \_gnd_net_\,
            in3 => \N__28582\,
            lcout => \elapsed_time_ns_1_RNIHG91B_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29584\,
            in2 => \_gnd_net_\,
            in3 => \N__29462\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28562\,
            in1 => \N__35190\,
            in2 => \_gnd_net_\,
            in3 => \N__32336\,
            lcout => \elapsed_time_ns_1_RNIVAQBB_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28976\,
            in1 => \N__35147\,
            in2 => \_gnd_net_\,
            in3 => \N__32337\,
            lcout => \elapsed_time_ns_1_RNI0CQBB_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_25_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28953\,
            in1 => \N__34514\,
            in2 => \_gnd_net_\,
            in3 => \N__32414\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49931\,
            ce => \N__28920\,
            sr => \N__49187\
        );

    \phase_controller_inst2.state_RNIG7JF_2_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28882\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28862\,
            lcout => \phase_controller_inst2.N_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__28702\,
            in1 => \N__28881\,
            in2 => \N__28868\,
            in3 => \N__29015\,
            lcout => \phase_controller_inst2.N_51_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29785\,
            in2 => \_gnd_net_\,
            in3 => \N__35994\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_165_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29935\,
            in2 => \_gnd_net_\,
            in3 => \N__29874\,
            lcout => \phase_controller_inst2.test_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_0_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__29086\,
            in1 => \N__28711\,
            in2 => \N__29072\,
            in3 => \N__29020\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49196\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110010101100"
        )
    port map (
            in0 => \N__28841\,
            in1 => \N__29087\,
            in2 => \N__28790\,
            in3 => \N__28748\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49196\
        );

    \phase_controller_inst2.state_1_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__28712\,
            in1 => \N__29019\,
            in2 => \_gnd_net_\,
            in3 => \N__28679\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49196\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__29786\,
            in1 => \N__35966\,
            in2 => \_gnd_net_\,
            in3 => \N__35996\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49196\
        );

    \phase_controller_inst2.start_timer_tr_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001101110011"
        )
    port map (
            in0 => \N__33351\,
            in1 => \N__29132\,
            in2 => \N__29117\,
            in3 => \N__29902\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49196\
        );

    \phase_controller_inst2.state_RNI9M3O_0_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29085\,
            in2 => \_gnd_net_\,
            in3 => \N__29068\,
            lcout => \phase_controller_inst2.N_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30928\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49906\,
            ce => 'H',
            sr => \N__49209\
        );

    \current_shift_inst.PI_CTRL.prop_term_29_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30784\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49903\,
            ce => 'H',
            sr => \N__49215\
        );

    \current_shift_inst.PI_CTRL.prop_term_30_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30757\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49903\,
            ce => 'H',
            sr => \N__49215\
        );

    \current_shift_inst.PI_CTRL.prop_term_28_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30808\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49903\,
            ce => 'H',
            sr => \N__49215\
        );

    \phase_controller_inst2.S2_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29021\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49222\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__31022\,
            in1 => \N__33207\,
            in2 => \N__31049\,
            in3 => \N__35814\,
            lcout => \phase_controller_inst1.N_49_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33934\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49993\,
            ce => \N__35099\,
            sr => \N__49129\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33865\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49993\,
            ce => \N__35099\,
            sr => \N__49129\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29200\,
            in1 => \N__29228\,
            in2 => \_gnd_net_\,
            in3 => \N__32165\,
            lcout => \elapsed_time_ns_1_RNIED91B_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29179\,
            in1 => \N__33830\,
            in2 => \_gnd_net_\,
            in3 => \N__32166\,
            lcout => \elapsed_time_ns_1_RNIGF91B_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34385\,
            in1 => \N__34458\,
            in2 => \N__34314\,
            in3 => \N__33465\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33537\,
            in2 => \_gnd_net_\,
            in3 => \N__33608\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33683\,
            in1 => \N__33758\,
            in2 => \N__29159\,
            in3 => \N__29156\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__35375\,
            in1 => \N__35440\,
            in2 => \_gnd_net_\,
            in3 => \N__29150\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__35150\,
            in1 => \N__29141\,
            in2 => \N__29135\,
            in3 => \N__30977\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__29416\,
            in1 => \_gnd_net_\,
            in2 => \N__29420\,
            in3 => \N__34640\,
            lcout => \elapsed_time_ns_1_RNI1CPBB_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29344\,
            in1 => \N__34045\,
            in2 => \_gnd_net_\,
            in3 => \N__32164\,
            lcout => \elapsed_time_ns_1_RNI3DOBB_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__29324\,
            in1 => \N__31579\,
            in2 => \N__29360\,
            in3 => \N__31556\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__31555\,
            in1 => \N__29323\,
            in2 => \N__31583\,
            in3 => \N__29356\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33969\,
            in1 => \N__32167\,
            in2 => \_gnd_net_\,
            in3 => \N__29374\,
            lcout => \elapsed_time_ns_1_RNI4EOBB_0_17\,
            ltout => \elapsed_time_ns_1_RNI4EOBB_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32169\,
            in1 => \_gnd_net_\,
            in2 => \N__29363\,
            in3 => \N__33970\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49974\,
            ce => \N__32703\,
            sr => \N__49141\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32168\,
            in1 => \N__29340\,
            in2 => \_gnd_net_\,
            in3 => \N__34046\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49974\,
            ce => \N__32703\,
            sr => \N__49141\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29314\,
            in1 => \N__32170\,
            in2 => \_gnd_net_\,
            in3 => \N__34243\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49974\,
            ce => \N__32703\,
            sr => \N__49141\
        );

    \phase_controller_inst1.start_timer_tr_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101011101"
        )
    port map (
            in0 => \N__29282\,
            in1 => \N__29454\,
            in2 => \N__33374\,
            in3 => \N__31979\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49967\,
            ce => 'H',
            sr => \N__49148\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__29453\,
            in1 => \N__29470\,
            in2 => \_gnd_net_\,
            in3 => \N__29571\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => \phase_controller_inst1.stoper_tr.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000111010"
        )
    port map (
            in0 => \N__29471\,
            in1 => \N__29577\,
            in2 => \N__29474\,
            in3 => \N__29548\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49967\,
            ce => 'H',
            sr => \N__49148\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29455\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49967\,
            ce => 'H',
            sr => \N__49148\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29570\,
            in2 => \_gnd_net_\,
            in3 => \N__29544\,
            lcout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29438\,
            in3 => \N__31218\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29749\,
            in1 => \N__33927\,
            in2 => \_gnd_net_\,
            in3 => \N__29435\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__49960\,
            ce => \N__29857\,
            sr => \N__49154\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29745\,
            in1 => \N__33864\,
            in2 => \_gnd_net_\,
            in3 => \N__29432\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__49960\,
            ce => \N__29857\,
            sr => \N__49154\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29750\,
            in1 => \N__33784\,
            in2 => \_gnd_net_\,
            in3 => \N__29429\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__49960\,
            ce => \N__29857\,
            sr => \N__49154\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29746\,
            in1 => \N__33705\,
            in2 => \_gnd_net_\,
            in3 => \N__29426\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__49960\,
            ce => \N__29857\,
            sr => \N__49154\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29751\,
            in1 => \N__33633\,
            in2 => \_gnd_net_\,
            in3 => \N__29423\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__49960\,
            ce => \N__29857\,
            sr => \N__49154\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29747\,
            in1 => \N__33561\,
            in2 => \_gnd_net_\,
            in3 => \N__29501\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__49960\,
            ce => \N__29857\,
            sr => \N__49154\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29752\,
            in1 => \N__33490\,
            in2 => \_gnd_net_\,
            in3 => \N__29498\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__49960\,
            ce => \N__29857\,
            sr => \N__49154\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29748\,
            in1 => \N__33417\,
            in2 => \_gnd_net_\,
            in3 => \N__29495\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__49960\,
            ce => \N__29857\,
            sr => \N__49154\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29709\,
            in1 => \N__34428\,
            in2 => \_gnd_net_\,
            in3 => \N__29492\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__49951\,
            ce => \N__29858\,
            sr => \N__49160\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29738\,
            in1 => \N__34347\,
            in2 => \_gnd_net_\,
            in3 => \N__29489\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__49951\,
            ce => \N__29858\,
            sr => \N__49160\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29706\,
            in1 => \N__34260\,
            in2 => \_gnd_net_\,
            in3 => \N__29486\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__49951\,
            ce => \N__29858\,
            sr => \N__49160\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29735\,
            in1 => \N__34191\,
            in2 => \_gnd_net_\,
            in3 => \N__29483\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__49951\,
            ce => \N__29858\,
            sr => \N__49160\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29707\,
            in1 => \N__34122\,
            in2 => \_gnd_net_\,
            in3 => \N__29480\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__49951\,
            ce => \N__29858\,
            sr => \N__49160\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29736\,
            in1 => \N__34062\,
            in2 => \_gnd_net_\,
            in3 => \N__29477\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__49951\,
            ce => \N__29858\,
            sr => \N__49160\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29708\,
            in1 => \N__33990\,
            in2 => \_gnd_net_\,
            in3 => \N__29528\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__49951\,
            ce => \N__29858\,
            sr => \N__49160\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29737\,
            in1 => \N__35029\,
            in2 => \_gnd_net_\,
            in3 => \N__29525\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__49951\,
            ce => \N__29858\,
            sr => \N__49160\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29731\,
            in1 => \N__34965\,
            in2 => \_gnd_net_\,
            in3 => \N__29522\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__49944\,
            ce => \N__29856\,
            sr => \N__49166\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29762\,
            in1 => \N__34878\,
            in2 => \_gnd_net_\,
            in3 => \N__29519\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__49944\,
            ce => \N__29856\,
            sr => \N__49166\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29732\,
            in1 => \N__34800\,
            in2 => \_gnd_net_\,
            in3 => \N__29516\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__49944\,
            ce => \N__29856\,
            sr => \N__49166\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29763\,
            in1 => \N__34734\,
            in2 => \_gnd_net_\,
            in3 => \N__29513\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__49944\,
            ce => \N__29856\,
            sr => \N__49166\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29733\,
            in1 => \N__34662\,
            in2 => \_gnd_net_\,
            in3 => \N__29510\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__49944\,
            ce => \N__29856\,
            sr => \N__49166\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29764\,
            in1 => \N__34591\,
            in2 => \_gnd_net_\,
            in3 => \N__29507\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__49944\,
            ce => \N__29856\,
            sr => \N__49166\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29734\,
            in1 => \N__34528\,
            in2 => \_gnd_net_\,
            in3 => \N__29504\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__49944\,
            ce => \N__29856\,
            sr => \N__49166\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29765\,
            in1 => \N__35545\,
            in2 => \_gnd_net_\,
            in3 => \N__29606\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__49944\,
            ce => \N__29856\,
            sr => \N__49166\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29739\,
            in1 => \N__35463\,
            in2 => \_gnd_net_\,
            in3 => \N__29603\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__49939\,
            ce => \N__29852\,
            sr => \N__49171\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29743\,
            in1 => \N__35391\,
            in2 => \_gnd_net_\,
            in3 => \N__29600\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__49939\,
            ce => \N__29852\,
            sr => \N__49171\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29740\,
            in1 => \N__35292\,
            in2 => \_gnd_net_\,
            in3 => \N__29597\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__49939\,
            ce => \N__29852\,
            sr => \N__49171\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29744\,
            in1 => \N__35206\,
            in2 => \_gnd_net_\,
            in3 => \N__29594\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__49939\,
            ce => \N__29852\,
            sr => \N__49171\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29741\,
            in1 => \N__35317\,
            in2 => \_gnd_net_\,
            in3 => \N__29591\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__49939\,
            ce => \N__29852\,
            sr => \N__49171\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__35233\,
            in1 => \N__29742\,
            in2 => \_gnd_net_\,
            in3 => \N__29588\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49939\,
            ce => \N__29852\,
            sr => \N__49171\
        );

    \phase_controller_inst1.state_0_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__33211\,
            in1 => \N__30020\,
            in2 => \N__30038\,
            in3 => \N__35825\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49932\,
            ce => 'H',
            sr => \N__49175\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110010101100"
        )
    port map (
            in0 => \N__29585\,
            in1 => \N__30037\,
            in2 => \N__31234\,
            in3 => \N__29552\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49932\,
            ce => 'H',
            sr => \N__49175\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30033\,
            in2 => \_gnd_net_\,
            in3 => \N__30019\,
            lcout => \phase_controller_inst1.N_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNILR64_4_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29994\,
            in2 => \_gnd_net_\,
            in3 => \N__33363\,
            lcout => \phase_controller_inst1_N_54\,
            ltout => \phase_controller_inst1_N_54_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_3_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__29880\,
            in1 => \N__29942\,
            in2 => \N__29909\,
            in3 => \N__29906\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49926\,
            ce => 'H',
            sr => \N__49181\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__29784\,
            in1 => \N__35965\,
            in2 => \_gnd_net_\,
            in3 => \N__35995\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_166_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__29812\,
            in1 => \N__31912\,
            in2 => \_gnd_net_\,
            in3 => \N__31950\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29783\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__37016\,
            in1 => \N__38579\,
            in2 => \_gnd_net_\,
            in3 => \N__41802\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38516\,
            in1 => \N__36953\,
            in2 => \_gnd_net_\,
            in3 => \N__41800\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => \current_shift_inst.control_input_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29639\,
            in3 => \N__32935\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49914\,
            ce => 'H',
            sr => \N__49192\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41801\,
            lcout => \current_shift_inst.N_1271_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__41803\,
            in1 => \N__38564\,
            in2 => \_gnd_net_\,
            in3 => \N__37001\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32915\,
            in1 => \N__30212\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32906\,
            in2 => \_gnd_net_\,
            in3 => \N__30173\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49197\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32894\,
            in3 => \N__30140\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49197\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32879\,
            in2 => \_gnd_net_\,
            in3 => \N__30110\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49197\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32867\,
            in2 => \_gnd_net_\,
            in3 => \N__30074\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49197\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32855\,
            in3 => \N__30041\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49197\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32840\,
            in2 => \_gnd_net_\,
            in3 => \N__30455\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49197\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32828\,
            in3 => \N__30425\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49197\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32807\,
            in3 => \N__30392\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_11_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49202\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33056\,
            in2 => \_gnd_net_\,
            in3 => \N__30362\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49202\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33044\,
            in3 => \N__30332\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49202\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33029\,
            in2 => \_gnd_net_\,
            in3 => \N__30302\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49202\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33017\,
            in2 => \_gnd_net_\,
            in3 => \N__30278\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49202\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33005\,
            in3 => \N__30245\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49202\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32990\,
            in2 => \_gnd_net_\,
            in3 => \N__30215\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49202\
        );

    \current_shift_inst.PI_CTRL.error_control_15_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32978\,
            in3 => \N__30701\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49202\
        );

    \current_shift_inst.PI_CTRL.error_control_16_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32963\,
            in3 => \N__30665\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_16\,
            ltout => OPEN,
            carryin => \bfn_11_21_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49205\
        );

    \current_shift_inst.PI_CTRL.error_control_17_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33173\,
            in2 => \_gnd_net_\,
            in3 => \N__30635\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49205\
        );

    \current_shift_inst.PI_CTRL.error_control_18_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33161\,
            in3 => \N__30602\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49205\
        );

    \current_shift_inst.PI_CTRL.error_control_19_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33146\,
            in2 => \_gnd_net_\,
            in3 => \N__30572\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49205\
        );

    \current_shift_inst.PI_CTRL.error_control_20_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33134\,
            in2 => \_gnd_net_\,
            in3 => \N__30545\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49205\
        );

    \current_shift_inst.PI_CTRL.error_control_21_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33122\,
            in3 => \N__30515\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49205\
        );

    \current_shift_inst.PI_CTRL.error_control_22_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33107\,
            in2 => \_gnd_net_\,
            in3 => \N__30491\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49205\
        );

    \current_shift_inst.PI_CTRL.error_control_23_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33095\,
            in3 => \N__30944\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49205\
        );

    \current_shift_inst.PI_CTRL.error_control_24_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33080\,
            in3 => \N__30914\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_24\,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49210\
        );

    \current_shift_inst.PI_CTRL.error_control_25_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33314\,
            in2 => \_gnd_net_\,
            in3 => \N__30884\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49210\
        );

    \current_shift_inst.PI_CTRL.error_control_26_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33302\,
            in3 => \N__30851\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49210\
        );

    \current_shift_inst.PI_CTRL.error_control_27_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33287\,
            in2 => \_gnd_net_\,
            in3 => \N__30824\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49210\
        );

    \current_shift_inst.PI_CTRL.error_control_28_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33275\,
            in2 => \_gnd_net_\,
            in3 => \N__30794\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49210\
        );

    \current_shift_inst.PI_CTRL.error_control_29_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33263\,
            in3 => \N__30767\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49210\
        );

    \current_shift_inst.PI_CTRL.error_control_30_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33230\,
            in2 => \_gnd_net_\,
            in3 => \N__30743\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_30\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49210\
        );

    \current_shift_inst.PI_CTRL.error_control_31_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__33245\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30740\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49210\
        );

    \phase_controller_inst1.stoper_hc.target_time_25_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44305\,
            in1 => \N__44276\,
            in2 => \_gnd_net_\,
            in3 => \N__50527\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50026\,
            ce => \N__49521\,
            sr => \N__49099\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50484\,
            in1 => \N__40248\,
            in2 => \_gnd_net_\,
            in3 => \N__43368\,
            lcout => \elapsed_time_ns_1_RNIV1DN9_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31071\,
            in1 => \N__34935\,
            in2 => \_gnd_net_\,
            in3 => \N__32324\,
            lcout => \elapsed_time_ns_1_RNI6GOBB_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_2_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__31047\,
            in1 => \N__35667\,
            in2 => \N__31028\,
            in3 => \N__35886\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49991\,
            ce => 'H',
            sr => \N__49115\
        );

    \phase_controller_inst1.state_RNIE87F_2_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31023\,
            in2 => \_gnd_net_\,
            in3 => \N__31046\,
            lcout => \phase_controller_inst1.N_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110010101100"
        )
    port map (
            in0 => \N__39551\,
            in1 => \N__31048\,
            in2 => \N__39455\,
            in3 => \N__39504\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49991\,
            ce => 'H',
            sr => \N__49115\
        );

    \phase_controller_inst1.test22_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__31027\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30988\,
            lcout => test22_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49991\,
            ce => 'H',
            sr => \N__49115\
        );

    \phase_controller_inst1.stoper_hc.target_time_21_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50493\,
            in1 => \N__40249\,
            in2 => \_gnd_net_\,
            in3 => \N__43369\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49983\,
            ce => \N__49465\,
            sr => \N__49123\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31247\,
            in1 => \N__31178\,
            in2 => \N__31256\,
            in3 => \N__31241\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_21_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31305\,
            in1 => \N__34777\,
            in2 => \_gnd_net_\,
            in3 => \N__32189\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49973\,
            ce => \N__32725\,
            sr => \N__49130\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35275\,
            in1 => \N__35189\,
            in2 => \N__35526\,
            in3 => \N__34512\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34706\,
            in1 => \N__34565\,
            in2 => \N__34644\,
            in3 => \N__34766\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34100\,
            in1 => \N__34029\,
            in2 => \N__34173\,
            in3 => \N__34229\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31217\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31189\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34830\,
            in1 => \N__34998\,
            in2 => \N__34934\,
            in3 => \N__33960\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31171\,
            in2 => \N__31136\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32704\,
            in1 => \N__31123\,
            in2 => \_gnd_net_\,
            in3 => \N__31109\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__49958\,
            ce => 'H',
            sr => \N__49142\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__32722\,
            in1 => \N__31106\,
            in2 => \N__31099\,
            in3 => \N__31079\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__49958\,
            ce => 'H',
            sr => \N__49142\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32705\,
            in1 => \N__31474\,
            in2 => \_gnd_net_\,
            in3 => \N__31460\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__49958\,
            ce => 'H',
            sr => \N__49142\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32723\,
            in1 => \N__31453\,
            in2 => \_gnd_net_\,
            in3 => \N__31439\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__49958\,
            ce => 'H',
            sr => \N__49142\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32706\,
            in1 => \N__31432\,
            in2 => \_gnd_net_\,
            in3 => \N__31418\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__49958\,
            ce => 'H',
            sr => \N__49142\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32724\,
            in1 => \N__31411\,
            in2 => \_gnd_net_\,
            in3 => \N__31397\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__49958\,
            ce => 'H',
            sr => \N__49142\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32707\,
            in1 => \N__31390\,
            in2 => \_gnd_net_\,
            in3 => \N__31376\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__49958\,
            ce => 'H',
            sr => \N__49142\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32715\,
            in1 => \N__31369\,
            in2 => \_gnd_net_\,
            in3 => \N__31355\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49149\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32708\,
            in1 => \N__31348\,
            in2 => \_gnd_net_\,
            in3 => \N__31334\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49149\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32712\,
            in1 => \N__31327\,
            in2 => \_gnd_net_\,
            in3 => \N__31313\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49149\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32709\,
            in1 => \N__31663\,
            in2 => \_gnd_net_\,
            in3 => \N__31649\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49149\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32713\,
            in1 => \N__31642\,
            in2 => \_gnd_net_\,
            in3 => \N__31628\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49149\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32710\,
            in1 => \N__31621\,
            in2 => \_gnd_net_\,
            in3 => \N__31607\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49149\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32714\,
            in1 => \N__31600\,
            in2 => \_gnd_net_\,
            in3 => \N__31586\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49149\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32711\,
            in1 => \N__31573\,
            in2 => \_gnd_net_\,
            in3 => \N__31559\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49149\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32689\,
            in1 => \N__31554\,
            in2 => \_gnd_net_\,
            in3 => \N__31538\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32672\,
            in1 => \N__31525\,
            in2 => \_gnd_net_\,
            in3 => \N__31511\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32690\,
            in1 => \N__31495\,
            in2 => \_gnd_net_\,
            in3 => \N__31481\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32673\,
            in1 => \N__31896\,
            in2 => \_gnd_net_\,
            in3 => \N__31874\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32691\,
            in1 => \N__31866\,
            in2 => \_gnd_net_\,
            in3 => \N__31847\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32674\,
            in1 => \N__31837\,
            in2 => \_gnd_net_\,
            in3 => \N__31823\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32692\,
            in1 => \N__31806\,
            in2 => \_gnd_net_\,
            in3 => \N__31790\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32675\,
            in1 => \N__31779\,
            in2 => \_gnd_net_\,
            in3 => \N__31763\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32665\,
            in1 => \N__31753\,
            in2 => \_gnd_net_\,
            in3 => \N__31739\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49161\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32669\,
            in1 => \N__31731\,
            in2 => \_gnd_net_\,
            in3 => \N__31715\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49161\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32666\,
            in1 => \N__31710\,
            in2 => \_gnd_net_\,
            in3 => \N__31694\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49161\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32670\,
            in1 => \N__31686\,
            in2 => \_gnd_net_\,
            in3 => \N__31670\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49161\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32667\,
            in1 => \N__32790\,
            in2 => \_gnd_net_\,
            in3 => \N__32774\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49161\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32671\,
            in1 => \N__32760\,
            in2 => \_gnd_net_\,
            in3 => \N__32741\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49161\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32668\,
            in1 => \N__32472\,
            in2 => \_gnd_net_\,
            in3 => \N__32477\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49161\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32448\,
            in1 => \N__34566\,
            in2 => \_gnd_net_\,
            in3 => \N__32413\,
            lcout => \elapsed_time_ns_1_RNI2DPBB_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34166\,
            in1 => \N__32001\,
            in2 => \_gnd_net_\,
            in3 => \N__32412\,
            lcout => \elapsed_time_ns_1_RNI1BOBB_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_3_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__31975\,
            in1 => \N__35678\,
            in2 => \N__35887\,
            in3 => \N__31964\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49919\,
            ce => 'H',
            sr => \N__49176\
        );

    \phase_controller_inst2.stoper_hc.running_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000101110"
        )
    port map (
            in0 => \N__31913\,
            in1 => \N__36682\,
            in2 => \N__31958\,
            in3 => \N__38391\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49919\,
            ce => 'H',
            sr => \N__49176\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111001001110"
        )
    port map (
            in0 => \N__35704\,
            in1 => \N__36128\,
            in2 => \N__36164\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49919\,
            ce => 'H',
            sr => \N__49176\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32948\,
            in2 => \N__32942\,
            in3 => \N__32934\,
            lcout => \current_shift_inst.control_input_1\,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35582\,
            in2 => \_gnd_net_\,
            in3 => \N__32897\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35576\,
            in2 => \_gnd_net_\,
            in3 => \N__32882\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35570\,
            in2 => \_gnd_net_\,
            in3 => \N__32870\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35564\,
            in2 => \_gnd_net_\,
            in3 => \N__32858\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35765\,
            in2 => \_gnd_net_\,
            in3 => \N__32843\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35759\,
            in2 => \_gnd_net_\,
            in3 => \N__32831\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35711\,
            in2 => \_gnd_net_\,
            in3 => \N__32816\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32813\,
            in2 => \_gnd_net_\,
            in3 => \N__32795\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33065\,
            in3 => \N__33047\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35594\,
            in2 => \_gnd_net_\,
            in3 => \N__33032\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38867\,
            in2 => \_gnd_net_\,
            in3 => \N__33020\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38894\,
            in2 => \_gnd_net_\,
            in3 => \N__33008\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39059\,
            in2 => \_gnd_net_\,
            in3 => \N__32993\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_12\,
            carryout => \current_shift_inst.control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39032\,
            in2 => \_gnd_net_\,
            in3 => \N__32981\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_13\,
            carryout => \current_shift_inst.control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39008\,
            in2 => \_gnd_net_\,
            in3 => \N__32966\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_14\,
            carryout => \current_shift_inst.control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35588\,
            in2 => \_gnd_net_\,
            in3 => \N__32951\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => \current_shift_inst.control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35747\,
            in2 => \_gnd_net_\,
            in3 => \N__33164\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_16\,
            carryout => \current_shift_inst.control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35753\,
            in2 => \_gnd_net_\,
            in3 => \N__33149\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_17\,
            carryout => \current_shift_inst.control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37232\,
            in2 => \_gnd_net_\,
            in3 => \N__33137\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_18\,
            carryout => \current_shift_inst.control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35741\,
            in2 => \_gnd_net_\,
            in3 => \N__33125\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_19\,
            carryout => \current_shift_inst.control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35735\,
            in2 => \_gnd_net_\,
            in3 => \N__33110\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_20\,
            carryout => \current_shift_inst.control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35729\,
            in2 => \_gnd_net_\,
            in3 => \N__33098\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_21\,
            carryout => \current_shift_inst.control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39152\,
            in2 => \_gnd_net_\,
            in3 => \N__33083\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_22\,
            carryout => \current_shift_inst.control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38843\,
            in2 => \_gnd_net_\,
            in3 => \N__33068\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \current_shift_inst.control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36008\,
            in2 => \_gnd_net_\,
            in3 => \N__33305\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_24\,
            carryout => \current_shift_inst.control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35717\,
            in2 => \_gnd_net_\,
            in3 => \N__33290\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_25\,
            carryout => \current_shift_inst.control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35723\,
            in2 => \_gnd_net_\,
            in3 => \N__33278\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_26\,
            carryout => \current_shift_inst.control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37145\,
            in2 => \_gnd_net_\,
            in3 => \N__33266\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_27\,
            carryout => \current_shift_inst.control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36002\,
            in2 => \_gnd_net_\,
            in3 => \N__33251\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_28\,
            carryout => \current_shift_inst.control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41873\,
            in2 => \_gnd_net_\,
            in3 => \N__33248\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33241\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__49268\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pll_inst.red_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_1_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__33386\,
            in1 => \N__33212\,
            in2 => \_gnd_net_\,
            in3 => \N__35798\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50028\,
            ce => 'H',
            sr => \N__49100\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__39450\,
            in1 => \N__39476\,
            in2 => \N__37345\,
            in3 => \N__49429\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50028\,
            ce => 'H',
            sr => \N__49100\
        );

    \phase_controller_inst1.stoper_hc.running_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011111100001100"
        )
    port map (
            in0 => \N__39505\,
            in1 => \N__39451\,
            in2 => \N__39549\,
            in3 => \N__39271\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50028\,
            ce => 'H',
            sr => \N__49100\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39251\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50028\,
            ce => 'H',
            sr => \N__49100\
        );

    \phase_controller_inst1.start_timer_hc_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__33395\,
            in1 => \N__33385\,
            in2 => \N__39257\,
            in3 => \N__33370\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50028\,
            ce => 'H',
            sr => \N__49100\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39228\,
            in1 => \N__42671\,
            in2 => \_gnd_net_\,
            in3 => \N__50496\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50015\,
            ce => \N__49543\,
            sr => \N__49105\
        );

    \phase_controller_inst1.stoper_hc.target_time_24_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44387\,
            in1 => \N__44340\,
            in2 => \_gnd_net_\,
            in3 => \N__50495\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50015\,
            ce => \N__49543\,
            sr => \N__49105\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50494\,
            in1 => \N__37937\,
            in2 => \_gnd_net_\,
            in3 => \N__42389\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50015\,
            ce => \N__49543\,
            sr => \N__49105\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42524\,
            in1 => \N__37912\,
            in2 => \_gnd_net_\,
            in3 => \N__50497\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50015\,
            ce => \N__49543\,
            sr => \N__49105\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__36316\,
            in1 => \N__37799\,
            in2 => \N__36344\,
            in3 => \N__37826\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50481\,
            in1 => \N__44341\,
            in2 => \_gnd_net_\,
            in3 => \N__44386\,
            lcout => \elapsed_time_ns_1_RNI25DN9_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42573\,
            in1 => \N__37948\,
            in2 => \_gnd_net_\,
            in3 => \N__50482\,
            lcout => \elapsed_time_ns_1_RNIH33T9_0_5\,
            ltout => \elapsed_time_ns_1_RNIH33T9_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50483\,
            in1 => \_gnd_net_\,
            in2 => \N__33401\,
            in3 => \N__42574\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50005\,
            ce => \N__49500\,
            sr => \N__49110\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44298\,
            in1 => \N__44272\,
            in2 => \_gnd_net_\,
            in3 => \N__50480\,
            lcout => \elapsed_time_ns_1_RNI36DN9_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__36383\,
            in1 => \N__37856\,
            in2 => \N__37613\,
            in3 => \N__36371\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50485\,
            in1 => \N__40276\,
            in2 => \_gnd_net_\,
            in3 => \N__43425\,
            lcout => \elapsed_time_ns_1_RNIU0DN9_0_20\,
            ltout => \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_20_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__43426\,
            in1 => \_gnd_net_\,
            in2 => \N__33398\,
            in3 => \N__50486\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49994\,
            ce => \N__49577\,
            sr => \N__49116\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36459\,
            in1 => \N__43555\,
            in2 => \_gnd_net_\,
            in3 => \N__50522\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49984\,
            ce => \N__49549\,
            sr => \N__49124\
        );

    \phase_controller_inst1.stoper_hc.target_time_27_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43985\,
            in1 => \N__37872\,
            in2 => \_gnd_net_\,
            in3 => \N__50523\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49984\,
            ce => \N__49549\,
            sr => \N__49124\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37936\,
            in1 => \N__42388\,
            in2 => \_gnd_net_\,
            in3 => \N__50526\,
            lcout => \elapsed_time_ns_1_RNIK63T9_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35663\,
            in2 => \_gnd_net_\,
            in3 => \N__35888\,
            lcout => \phase_controller_inst1.test_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33790\,
            in2 => \N__33938\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__49968\,
            ce => \N__35105\,
            sr => \N__49137\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33712\,
            in2 => \N__33869\,
            in3 => \N__33794\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__49968\,
            ce => \N__35105\,
            sr => \N__49137\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33791\,
            in2 => \N__33644\,
            in3 => \N__33719\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__49968\,
            ce => \N__35105\,
            sr => \N__49137\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33568\,
            in2 => \N__33716\,
            in3 => \N__33647\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__49968\,
            ce => \N__35105\,
            sr => \N__49137\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33643\,
            in2 => \N__33502\,
            in3 => \N__33575\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__49968\,
            ce => \N__35105\,
            sr => \N__49137\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33424\,
            in2 => \N__33572\,
            in3 => \N__33506\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__49968\,
            ce => \N__35105\,
            sr => \N__49137\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34429\,
            in2 => \N__33503\,
            in3 => \N__33431\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__49968\,
            ce => \N__35105\,
            sr => \N__49137\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34348\,
            in2 => \N__33428\,
            in3 => \N__34439\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__49968\,
            ce => \N__35105\,
            sr => \N__49137\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34267\,
            in2 => \N__34436\,
            in3 => \N__34355\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__49961\,
            ce => \N__35104\,
            sr => \N__49143\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34198\,
            in2 => \N__34352\,
            in3 => \N__34274\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__49961\,
            ce => \N__35104\,
            sr => \N__49143\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34129\,
            in2 => \N__34271\,
            in3 => \N__34205\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__49961\,
            ce => \N__35104\,
            sr => \N__49143\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34069\,
            in2 => \N__34202\,
            in3 => \N__34136\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__49961\,
            ce => \N__35104\,
            sr => \N__49143\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33997\,
            in2 => \N__34133\,
            in3 => \N__34076\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__49961\,
            ce => \N__35104\,
            sr => \N__49143\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35035\,
            in2 => \N__34073\,
            in3 => \N__34004\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__49961\,
            ce => \N__35104\,
            sr => \N__49143\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34972\,
            in2 => \N__34001\,
            in3 => \N__33941\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__49961\,
            ce => \N__35104\,
            sr => \N__49143\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35036\,
            in2 => \N__34891\,
            in3 => \N__34982\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__49961\,
            ce => \N__35104\,
            sr => \N__49143\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34807\,
            in2 => \N__34979\,
            in3 => \N__34895\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__49952\,
            ce => \N__35100\,
            sr => \N__49150\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34741\,
            in2 => \N__34892\,
            in3 => \N__34814\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__49952\,
            ce => \N__35100\,
            sr => \N__49150\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34669\,
            in2 => \N__34811\,
            in3 => \N__34748\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__49952\,
            ce => \N__35100\,
            sr => \N__49150\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34597\,
            in2 => \N__34745\,
            in3 => \N__34676\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__49952\,
            ce => \N__35100\,
            sr => \N__49150\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34534\,
            in2 => \N__34673\,
            in3 => \N__34601\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__49952\,
            ce => \N__35100\,
            sr => \N__49150\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34598\,
            in2 => \N__35557\,
            in3 => \N__34538\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__49952\,
            ce => \N__35100\,
            sr => \N__49150\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34535\,
            in2 => \N__35480\,
            in3 => \N__34472\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__49952\,
            ce => \N__35100\,
            sr => \N__49150\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35398\,
            in2 => \N__35558\,
            in3 => \N__35483\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__49952\,
            ce => \N__35100\,
            sr => \N__49150\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35299\,
            in2 => \N__35479\,
            in3 => \N__35402\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__49945\,
            ce => \N__35086\,
            sr => \N__49156\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35399\,
            in2 => \N__35218\,
            in3 => \N__35324\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__49945\,
            ce => \N__35086\,
            sr => \N__49156\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35321\,
            in2 => \N__35303\,
            in3 => \N__35240\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__49945\,
            ce => \N__35086\,
            sr => \N__49156\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35237\,
            in2 => \N__35219\,
            in3 => \N__35156\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__49945\,
            ce => \N__35086\,
            sr => \N__49156\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35153\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => \N__35086\,
            sr => \N__49156\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35705\,
            in2 => \_gnd_net_\,
            in3 => \N__36156\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_163_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__36157\,
            in1 => \N__35700\,
            in2 => \_gnd_net_\,
            in3 => \N__36124\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_164_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38594\,
            in1 => \N__37025\,
            in2 => \_gnd_net_\,
            in3 => \N__41837\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35699\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.test_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__35671\,
            in1 => \N__35605\,
            in2 => \_gnd_net_\,
            in3 => \N__35874\,
            lcout => test_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49921\,
            ce => 'H',
            sr => \N__49177\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38549\,
            in1 => \N__36986\,
            in2 => \_gnd_net_\,
            in3 => \N__41810\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__41811\,
            in1 => \_gnd_net_\,
            in2 => \N__38735\,
            in3 => \N__37115\,
            lcout => \current_shift_inst.control_input_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__36938\,
            in1 => \N__38498\,
            in2 => \_gnd_net_\,
            in3 => \N__41804\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__41805\,
            in1 => \_gnd_net_\,
            in2 => \N__38480\,
            in3 => \N__36926\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38462\,
            in1 => \N__36911\,
            in2 => \_gnd_net_\,
            in3 => \N__41806\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__41807\,
            in1 => \N__38447\,
            in2 => \_gnd_net_\,
            in3 => \N__37064\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__37049\,
            in1 => \N__38624\,
            in2 => \_gnd_net_\,
            in3 => \N__41808\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__41809\,
            in1 => \N__38609\,
            in2 => \_gnd_net_\,
            in3 => \N__37037\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__41865\,
            in1 => \N__37094\,
            in2 => \_gnd_net_\,
            in3 => \N__38699\,
            lcout => \current_shift_inst.control_input_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001111"
        )
    port map (
            in0 => \N__37106\,
            in1 => \_gnd_net_\,
            in2 => \N__38717\,
            in3 => \N__41864\,
            lcout => \current_shift_inst.control_input_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__41866\,
            in1 => \_gnd_net_\,
            in2 => \N__38669\,
            in3 => \N__37076\,
            lcout => \current_shift_inst.control_input_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38651\,
            in1 => \N__37199\,
            in2 => \_gnd_net_\,
            in3 => \N__41867\,
            lcout => \current_shift_inst.control_input_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__41868\,
            in1 => \N__37190\,
            in2 => \_gnd_net_\,
            in3 => \N__38636\,
            lcout => \current_shift_inst.control_input_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38786\,
            in1 => \N__37157\,
            in2 => \_gnd_net_\,
            in3 => \N__41871\,
            lcout => \current_shift_inst.control_input_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__41870\,
            in1 => \N__38804\,
            in2 => \_gnd_net_\,
            in3 => \N__37166\,
            lcout => \current_shift_inst.control_input_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38822\,
            in1 => \N__37175\,
            in2 => \_gnd_net_\,
            in3 => \N__41869\,
            lcout => \current_shift_inst.control_input_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41872\,
            lcout => \current_shift_inst.control_input_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35957\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35933\,
            ce => 'H',
            sr => \N__49198\
        );

    \delay_measurement_inst.start_timer_tr_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35958\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35933\,
            ce => 'H',
            sr => \N__49198\
        );

    \current_shift_inst.stop_timer_s1_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__37463\,
            in1 => \N__35889\,
            in2 => \N__37421\,
            in3 => \N__35911\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49203\
        );

    \phase_controller_inst1.S1_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35890\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49203\
        );

    \current_shift_inst.start_timer_s1_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__35910\,
            in1 => \N__37461\,
            in2 => \_gnd_net_\,
            in3 => \N__35894\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49899\,
            ce => 'H',
            sr => \N__49206\
        );

    \current_shift_inst.timer_s1.running_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__37462\,
            in1 => \N__37416\,
            in2 => \_gnd_net_\,
            in3 => \N__37442\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49899\,
            ce => 'H',
            sr => \N__49206\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37420\,
            in2 => \_gnd_net_\,
            in3 => \N__37439\,
            lcout => \current_shift_inst.timer_s1.N_161_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_13_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35824\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49894\,
            ce => 'H',
            sr => \N__49232\
        );

    \delay_measurement_inst.stop_timer_hc_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36109\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36092\,
            ce => 'H',
            sr => \N__49091\
        );

    \delay_measurement_inst.start_timer_hc_LC_14_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36108\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36092\,
            ce => 'H',
            sr => \N__49091\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37335\,
            in1 => \N__37370\,
            in2 => \N__36083\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_14_4_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37382\,
            in2 => \N__36074\,
            in3 => \N__37319\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36065\,
            in2 => \N__36059\,
            in3 => \N__37300\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37376\,
            in2 => \N__36050\,
            in3 => \N__37582\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36041\,
            in2 => \N__36032\,
            in3 => \N__37567\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36014\,
            in2 => \N__36023\,
            in3 => \N__37552\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36245\,
            in2 => \N__37391\,
            in3 => \N__37537\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36239\,
            in2 => \N__36233\,
            in3 => \N__37522\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41108\,
            in2 => \N__36224\,
            in3 => \N__37507\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37492\,
            in1 => \N__41075\,
            in2 => \N__36215\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41039\,
            in2 => \N__36206\,
            in3 => \N__37477\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42683\,
            in2 => \N__36197\,
            in3 => \N__37723\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37708\,
            in1 => \N__39794\,
            in2 => \N__36185\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37693\,
            in1 => \N__40820\,
            in2 => \N__36176\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36470\,
            in2 => \N__36269\,
            in3 => \N__37678\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40913\,
            in2 => \N__40985\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36350\,
            in2 => \N__36281\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36356\,
            in2 => \N__36260\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39680\,
            in2 => \N__39635\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36251\,
            in2 => \N__36305\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36389\,
            in2 => \N__36407\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39356\,
            in2 => \N__39413\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39806\,
            in2 => \N__39590\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36410\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100010000"
        )
    port map (
            in0 => \N__37746\,
            in1 => \N__37764\,
            in2 => \N__37364\,
            in3 => \N__36398\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011101111"
        )
    port map (
            in0 => \N__36397\,
            in1 => \N__37363\,
            in2 => \N__37769\,
            in3 => \N__37747\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__36382\,
            in1 => \N__37851\,
            in2 => \N__37612\,
            in3 => \N__36370\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37876\,
            in1 => \N__43984\,
            in2 => \_gnd_net_\,
            in3 => \N__50500\,
            lcout => \elapsed_time_ns_1_RNI58DN9_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50499\,
            in1 => \N__42513\,
            in2 => \_gnd_net_\,
            in3 => \N__37911\,
            lcout => \elapsed_time_ns_1_RNII43T9_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__36296\,
            in1 => \N__37633\,
            in2 => \N__37658\,
            in3 => \N__36487\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101100001010"
        )
    port map (
            in0 => \N__36343\,
            in1 => \N__37821\,
            in2 => \N__37798\,
            in3 => \N__36320\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__36292\,
            in1 => \N__37653\,
            in2 => \N__36488\,
            in3 => \N__37632\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43554\,
            in1 => \N__36461\,
            in2 => \_gnd_net_\,
            in3 => \N__50394\,
            lcout => \elapsed_time_ns_1_RNI57CN9_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__43489\,
            in1 => \_gnd_net_\,
            in2 => \N__50498\,
            in3 => \N__36433\,
            lcout => \elapsed_time_ns_1_RNI68CN9_0_19\,
            ltout => \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43490\,
            in2 => \N__36491\,
            in3 => \N__50396\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49995\,
            ce => \N__49548\,
            sr => \N__49117\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42867\,
            in1 => \N__50390\,
            in2 => \_gnd_net_\,
            in3 => \N__37888\,
            lcout => \elapsed_time_ns_1_RNI24CN9_0_15\,
            ltout => \elapsed_time_ns_1_RNI24CN9_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50395\,
            in1 => \_gnd_net_\,
            in2 => \N__36473\,
            in3 => \N__42868\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49995\,
            ce => \N__49548\,
            sr => \N__49117\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__36614\,
            in1 => \N__36637\,
            in2 => \N__36422\,
            in3 => \N__36443\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__36442\,
            in1 => \N__36613\,
            in2 => \N__36641\,
            in3 => \N__36418\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36460\,
            in1 => \N__43559\,
            in2 => \_gnd_net_\,
            in3 => \N__50518\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49985\,
            ce => \N__45112\,
            sr => \N__49125\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50516\,
            in1 => \N__43488\,
            in2 => \_gnd_net_\,
            in3 => \N__36434\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49985\,
            ce => \N__45112\,
            sr => \N__49125\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39233\,
            in1 => \N__42670\,
            in2 => \_gnd_net_\,
            in3 => \N__50519\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49985\,
            ce => \N__45112\,
            sr => \N__49125\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50517\,
            in1 => \N__39299\,
            in2 => \_gnd_net_\,
            in3 => \N__42635\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49985\,
            ce => \N__45112\,
            sr => \N__49125\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36548\,
            in2 => \N__38162\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36874\,
            in1 => \N__38120\,
            in2 => \_gnd_net_\,
            in3 => \N__36530\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__49975\,
            ce => 'H',
            sr => \N__49131\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__36878\,
            in1 => \N__38089\,
            in2 => \N__36527\,
            in3 => \N__36506\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__49975\,
            ce => 'H',
            sr => \N__49131\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36875\,
            in1 => \N__38069\,
            in2 => \_gnd_net_\,
            in3 => \N__36503\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__49975\,
            ce => 'H',
            sr => \N__49131\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36879\,
            in1 => \N__38036\,
            in2 => \_gnd_net_\,
            in3 => \N__36500\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__49975\,
            ce => 'H',
            sr => \N__49131\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36876\,
            in1 => \N__38012\,
            in2 => \_gnd_net_\,
            in3 => \N__36497\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__49975\,
            ce => 'H',
            sr => \N__49131\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36880\,
            in1 => \N__37981\,
            in2 => \_gnd_net_\,
            in3 => \N__36494\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__49975\,
            ce => 'H',
            sr => \N__49131\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36877\,
            in1 => \N__38345\,
            in2 => \_gnd_net_\,
            in3 => \N__36575\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__49975\,
            ce => 'H',
            sr => \N__49131\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36866\,
            in1 => \N__38324\,
            in2 => \_gnd_net_\,
            in3 => \N__36572\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__49969\,
            ce => 'H',
            sr => \N__49138\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36831\,
            in1 => \N__38303\,
            in2 => \_gnd_net_\,
            in3 => \N__36569\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__49969\,
            ce => 'H',
            sr => \N__49138\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36863\,
            in1 => \N__38282\,
            in2 => \_gnd_net_\,
            in3 => \N__36566\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__49969\,
            ce => 'H',
            sr => \N__49138\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36832\,
            in1 => \N__38261\,
            in2 => \_gnd_net_\,
            in3 => \N__36563\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__49969\,
            ce => 'H',
            sr => \N__49138\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36864\,
            in1 => \N__38240\,
            in2 => \_gnd_net_\,
            in3 => \N__36560\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__49969\,
            ce => 'H',
            sr => \N__49138\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36833\,
            in1 => \N__38219\,
            in2 => \_gnd_net_\,
            in3 => \N__36557\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__49969\,
            ce => 'H',
            sr => \N__49138\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36865\,
            in1 => \N__38189\,
            in2 => \_gnd_net_\,
            in3 => \N__36554\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__49969\,
            ce => 'H',
            sr => \N__49138\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36834\,
            in1 => \N__39766\,
            in2 => \_gnd_net_\,
            in3 => \N__36551\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__49969\,
            ce => 'H',
            sr => \N__49138\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36851\,
            in1 => \N__39742\,
            in2 => \_gnd_net_\,
            in3 => \N__36644\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49144\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36855\,
            in1 => \N__36631\,
            in2 => \_gnd_net_\,
            in3 => \N__36617\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49144\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36852\,
            in1 => \N__36612\,
            in2 => \_gnd_net_\,
            in3 => \N__36596\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49144\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36856\,
            in1 => \N__40303\,
            in2 => \_gnd_net_\,
            in3 => \N__36593\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49144\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36853\,
            in1 => \N__40327\,
            in2 => \_gnd_net_\,
            in3 => \N__36590\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49144\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36857\,
            in1 => \N__40164\,
            in2 => \_gnd_net_\,
            in3 => \N__36587\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49144\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36854\,
            in1 => \N__40147\,
            in2 => \_gnd_net_\,
            in3 => \N__36584\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49144\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36858\,
            in1 => \N__44436\,
            in2 => \_gnd_net_\,
            in3 => \N__36581\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49144\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36859\,
            in1 => \N__44410\,
            in2 => \_gnd_net_\,
            in3 => \N__36578\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__49953\,
            ce => 'H',
            sr => \N__49151\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36867\,
            in1 => \N__40027\,
            in2 => \_gnd_net_\,
            in3 => \N__36899\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__49953\,
            ce => 'H',
            sr => \N__49151\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36860\,
            in1 => \N__40063\,
            in2 => \_gnd_net_\,
            in3 => \N__36896\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__49953\,
            ce => 'H',
            sr => \N__49151\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36868\,
            in1 => \N__39937\,
            in2 => \_gnd_net_\,
            in3 => \N__36893\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__49953\,
            ce => 'H',
            sr => \N__49151\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36861\,
            in1 => \N__39913\,
            in2 => \_gnd_net_\,
            in3 => \N__36890\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__49953\,
            ce => 'H',
            sr => \N__49151\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36869\,
            in1 => \N__44191\,
            in2 => \_gnd_net_\,
            in3 => \N__36887\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__49953\,
            ce => 'H',
            sr => \N__49151\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36862\,
            in1 => \N__44167\,
            in2 => \_gnd_net_\,
            in3 => \N__36884\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49953\,
            ce => 'H',
            sr => \N__49151\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__36870\,
            in1 => \N__36728\,
            in2 => \N__36701\,
            in3 => \N__38157\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49953\,
            ce => 'H',
            sr => \N__49151\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46375\,
            in1 => \N__45832\,
            in2 => \N__46880\,
            in3 => \N__40582\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47758\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49946\,
            ce => \N__47792\,
            sr => \N__49157\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46376\,
            in1 => \N__45833\,
            in2 => \N__46879\,
            in3 => \N__40583\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45831\,
            in1 => \N__46377\,
            in2 => \N__46930\,
            in3 => \N__40613\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44627\,
            in2 => \N__45653\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45023\,
            in1 => \N__40473\,
            in2 => \N__40505\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46252\,
            in2 => \N__36968\,
            in3 => \N__45024\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36959\,
            in2 => \N__46439\,
            in3 => \N__36941\,
            lcout => \current_shift_inst.un38_control_input_0_s0_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46256\,
            in2 => \N__41315\,
            in3 => \N__36929\,
            lcout => \current_shift_inst.un38_control_input_0_s0_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44525\,
            in2 => \N__46440\,
            in3 => \N__36914\,
            lcout => \current_shift_inst.un38_control_input_0_s0_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46260\,
            in2 => \N__38948\,
            in3 => \N__36902\,
            lcout => \current_shift_inst.un38_control_input_0_s0_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37133\,
            in2 => \N__46441\,
            in3 => \N__37052\,
            lcout => \current_shift_inst.un38_control_input_0_s0_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46280\,
            in2 => \N__46673\,
            in3 => \N__37040\,
            lcout => \current_shift_inst.un38_control_input_0_s0_8\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40559\,
            in2 => \N__46446\,
            in3 => \N__37028\,
            lcout => \current_shift_inst.un38_control_input_0_s0_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46284\,
            in2 => \N__46058\,
            in3 => \N__37019\,
            lcout => \current_shift_inst.un38_control_input_0_s0_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38753\,
            in2 => \N__46447\,
            in3 => \N__37004\,
            lcout => \current_shift_inst.un38_control_input_0_s0_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46288\,
            in2 => \N__41651\,
            in3 => \N__36989\,
            lcout => \current_shift_inst.un38_control_input_0_s0_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38747\,
            in2 => \N__46448\,
            in3 => \N__36977\,
            lcout => \current_shift_inst.un38_control_input_0_s0_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46292\,
            in2 => \N__38933\,
            in3 => \N__36974\,
            lcout => \current_shift_inst.un38_control_input_0_s0_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45179\,
            in2 => \N__46449\,
            in3 => \N__36971\,
            lcout => \current_shift_inst.un38_control_input_0_s0_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46450\,
            in2 => \N__41378\,
            in3 => \N__37124\,
            lcout => \current_shift_inst.un38_control_input_0_s0_16\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37217\,
            in2 => \N__46593\,
            in3 => \N__37121\,
            lcout => \current_shift_inst.un38_control_input_0_s0_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46454\,
            in2 => \N__37262\,
            in3 => \N__37118\,
            lcout => \current_shift_inst.un38_control_input_0_s0_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38999\,
            in2 => \N__46594\,
            in3 => \N__37109\,
            lcout => \current_shift_inst.un38_control_input_0_s0_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46458\,
            in2 => \N__37286\,
            in3 => \N__37097\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38993\,
            in2 => \N__46595\,
            in3 => \N__37082\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46462\,
            in2 => \N__37274\,
            in3 => \N__37079\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37250\,
            in2 => \N__46596\,
            in3 => \N__37067\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37223\,
            in2 => \N__46597\,
            in3 => \N__37193\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46469\,
            in2 => \N__39194\,
            in3 => \N__37184\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38954\,
            in2 => \N__46598\,
            in3 => \N__37181\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46473\,
            in2 => \N__39176\,
            in3 => \N__37178\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37208\,
            in2 => \N__46599\,
            in3 => \N__37169\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46477\,
            in2 => \N__39143\,
            in3 => \N__37160\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39332\,
            in2 => \N__46600\,
            in3 => \N__37151\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010100110101"
        )
    port map (
            in0 => \N__38768\,
            in1 => \N__40541\,
            in2 => \N__41863\,
            in3 => \N__37148\,
            lcout => \current_shift_inst.control_input_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45874\,
            in1 => \N__46561\,
            in2 => \N__47305\,
            in3 => \N__40708\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46564\,
            in1 => \N__45877\,
            in2 => \N__47474\,
            in3 => \N__45473\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45878\,
            in1 => \N__46562\,
            in2 => \N__42185\,
            in3 => \N__47383\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__46560\,
            in1 => \N__45876\,
            in2 => \N__41924\,
            in3 => \N__47554\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45879\,
            in1 => \N__46563\,
            in2 => \N__47345\,
            in3 => \N__45170\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38684\,
            in1 => \N__37241\,
            in2 => \_gnd_net_\,
            in3 => \N__41861\,
            lcout => \current_shift_inst.control_input_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45880\,
            in1 => \N__46565\,
            in2 => \N__48059\,
            in3 => \N__42056\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__46566\,
            in1 => \N__47599\,
            in2 => \N__45638\,
            in3 => \N__45875\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45955\,
            in1 => \N__47876\,
            in2 => \N__46651\,
            in3 => \N__41720\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37440\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__37460\,
            in1 => \N__37441\,
            in2 => \_gnd_net_\,
            in3 => \N__37415\,
            lcout => \current_shift_inst.timer_s1.N_162_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50477\,
            in1 => \N__40216\,
            in2 => \_gnd_net_\,
            in3 => \N__42455\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50042\,
            ce => \N__49565\,
            sr => \N__49092\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39567\,
            in1 => \N__43701\,
            in2 => \_gnd_net_\,
            in3 => \N__50479\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50042\,
            ce => \N__49565\,
            sr => \N__49092\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__39288\,
            in1 => \_gnd_net_\,
            in2 => \N__50525\,
            in3 => \N__42631\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50042\,
            ce => \N__49565\,
            sr => \N__49092\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44480\,
            in1 => \N__44516\,
            in2 => \_gnd_net_\,
            in3 => \N__50478\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50042\,
            ce => \N__49565\,
            sr => \N__49092\
        );

    \phase_controller_inst1.stoper_hc.target_time_26_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50473\,
            in1 => \N__39996\,
            in2 => \_gnd_net_\,
            in3 => \N__44063\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50042\,
            ce => \N__49565\,
            sr => \N__49092\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39419\,
            in2 => \N__37349\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_5_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49356\,
            in1 => \N__37318\,
            in2 => \_gnd_net_\,
            in3 => \N__37304\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__50036\,
            ce => 'H',
            sr => \N__49095\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__49387\,
            in1 => \N__37301\,
            in2 => \N__39206\,
            in3 => \N__37289\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__50036\,
            ce => 'H',
            sr => \N__49095\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49357\,
            in1 => \N__37583\,
            in2 => \_gnd_net_\,
            in3 => \N__37571\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__50036\,
            ce => 'H',
            sr => \N__49095\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49388\,
            in1 => \N__37568\,
            in2 => \_gnd_net_\,
            in3 => \N__37556\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__50036\,
            ce => 'H',
            sr => \N__49095\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49358\,
            in1 => \N__37553\,
            in2 => \_gnd_net_\,
            in3 => \N__37541\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__50036\,
            ce => 'H',
            sr => \N__49095\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49389\,
            in1 => \N__37538\,
            in2 => \_gnd_net_\,
            in3 => \N__37526\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__50036\,
            ce => 'H',
            sr => \N__49095\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49359\,
            in1 => \N__37523\,
            in2 => \_gnd_net_\,
            in3 => \N__37511\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__50036\,
            ce => 'H',
            sr => \N__49095\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49525\,
            in1 => \N__37508\,
            in2 => \_gnd_net_\,
            in3 => \N__37496\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_6_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__50029\,
            ce => 'H',
            sr => \N__49101\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49433\,
            in1 => \N__37493\,
            in2 => \_gnd_net_\,
            in3 => \N__37481\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__50029\,
            ce => 'H',
            sr => \N__49101\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49522\,
            in1 => \N__37478\,
            in2 => \_gnd_net_\,
            in3 => \N__37466\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__50029\,
            ce => 'H',
            sr => \N__49101\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49434\,
            in1 => \N__37724\,
            in2 => \_gnd_net_\,
            in3 => \N__37712\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__50029\,
            ce => 'H',
            sr => \N__49101\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49523\,
            in1 => \N__37709\,
            in2 => \_gnd_net_\,
            in3 => \N__37697\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__50029\,
            ce => 'H',
            sr => \N__49101\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49435\,
            in1 => \N__37694\,
            in2 => \_gnd_net_\,
            in3 => \N__37682\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__50029\,
            ce => 'H',
            sr => \N__49101\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49524\,
            in1 => \N__37679\,
            in2 => \_gnd_net_\,
            in3 => \N__37667\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__50029\,
            ce => 'H',
            sr => \N__49101\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49436\,
            in1 => \N__40927\,
            in2 => \_gnd_net_\,
            in3 => \N__37664\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__50029\,
            ce => 'H',
            sr => \N__49101\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49526\,
            in1 => \N__40953\,
            in2 => \_gnd_net_\,
            in3 => \N__37661\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__50016\,
            ce => 'H',
            sr => \N__49106\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49461\,
            in1 => \N__37657\,
            in2 => \_gnd_net_\,
            in3 => \N__37637\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__50016\,
            ce => 'H',
            sr => \N__49106\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49527\,
            in1 => \N__37634\,
            in2 => \_gnd_net_\,
            in3 => \N__37616\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__50016\,
            ce => 'H',
            sr => \N__49106\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49462\,
            in1 => \N__37608\,
            in2 => \_gnd_net_\,
            in3 => \N__37586\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__50016\,
            ce => 'H',
            sr => \N__49106\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49528\,
            in1 => \N__37855\,
            in2 => \_gnd_net_\,
            in3 => \N__37835\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__50016\,
            ce => 'H',
            sr => \N__49106\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49463\,
            in1 => \N__39652\,
            in2 => \_gnd_net_\,
            in3 => \N__37832\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__50016\,
            ce => 'H',
            sr => \N__49106\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49529\,
            in1 => \N__39668\,
            in2 => \_gnd_net_\,
            in3 => \N__37829\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__50016\,
            ce => 'H',
            sr => \N__49106\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49464\,
            in1 => \N__37822\,
            in2 => \_gnd_net_\,
            in3 => \N__37802\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__50016\,
            ce => 'H',
            sr => \N__49106\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49469\,
            in1 => \N__37794\,
            in2 => \_gnd_net_\,
            in3 => \N__37772\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__50006\,
            ce => 'H',
            sr => \N__49111\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49578\,
            in1 => \N__37768\,
            in2 => \_gnd_net_\,
            in3 => \N__37751\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__50006\,
            ce => 'H',
            sr => \N__49111\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49470\,
            in1 => \N__37748\,
            in2 => \_gnd_net_\,
            in3 => \N__37733\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__50006\,
            ce => 'H',
            sr => \N__49111\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49579\,
            in1 => \N__39370\,
            in2 => \_gnd_net_\,
            in3 => \N__37730\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__50006\,
            ce => 'H',
            sr => \N__49111\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49471\,
            in1 => \N__39396\,
            in2 => \_gnd_net_\,
            in3 => \N__37727\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__50006\,
            ce => 'H',
            sr => \N__49111\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49580\,
            in1 => \N__39821\,
            in2 => \_gnd_net_\,
            in3 => \N__37961\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__50006\,
            ce => 'H',
            sr => \N__49111\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49472\,
            in1 => \N__39836\,
            in2 => \_gnd_net_\,
            in3 => \N__37958\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50006\,
            ce => 'H',
            sr => \N__49111\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50330\,
            in1 => \N__42578\,
            in2 => \_gnd_net_\,
            in3 => \N__37955\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49996\,
            ce => \N__45115\,
            sr => \N__49118\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50331\,
            in1 => \N__37935\,
            in2 => \_gnd_net_\,
            in3 => \N__42384\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49996\,
            ce => \N__45115\,
            sr => \N__49118\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37913\,
            in1 => \N__42520\,
            in2 => \_gnd_net_\,
            in3 => \N__50333\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49996\,
            ce => \N__45115\,
            sr => \N__49118\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50328\,
            in1 => \N__44473\,
            in2 => \_gnd_net_\,
            in3 => \N__44512\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49996\,
            ce => \N__45115\,
            sr => \N__49118\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42872\,
            in1 => \N__50332\,
            in2 => \_gnd_net_\,
            in3 => \N__37889\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49996\,
            ce => \N__45115\,
            sr => \N__49118\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50329\,
            in1 => \N__39575\,
            in2 => \_gnd_net_\,
            in3 => \N__43703\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49996\,
            ce => \N__45115\,
            sr => \N__49118\
        );

    \phase_controller_inst2.stoper_hc.target_time_27_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50520\,
            in1 => \N__37877\,
            in2 => \_gnd_net_\,
            in3 => \N__43983\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49996\,
            ce => \N__45115\,
            sr => \N__49118\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38132\,
            in2 => \N__38171\,
            in3 => \N__38161\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38126\,
            in2 => \N__38108\,
            in3 => \N__38119\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38075\,
            in2 => \N__38099\,
            in3 => \N__38090\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38068\,
            in1 => \N__38057\,
            in2 => \N__38051\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38042\,
            in2 => \N__38024\,
            in3 => \N__38035\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38011\,
            in1 => \N__38000\,
            in2 => \N__37994\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37982\,
            in1 => \N__37967\,
            in2 => \N__40193\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38351\,
            in2 => \N__38333\,
            in3 => \N__38344\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40184\,
            in2 => \N__38312\,
            in3 => \N__38323\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40391\,
            in2 => \N__38291\,
            in3 => \N__38302\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40397\,
            in2 => \N__38270\,
            in3 => \N__38281\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40385\,
            in2 => \N__38249\,
            in3 => \N__38260\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41228\,
            in2 => \N__38228\,
            in3 => \N__38239\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38218\,
            in1 => \N__38207\,
            in2 => \N__40094\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38177\,
            in2 => \N__38201\,
            in3 => \N__38188\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39782\,
            in2 => \N__39728\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38429\,
            in2 => \N__38417\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40289\,
            in2 => \N__40343\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40127\,
            in2 => \N__40178\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44396\,
            in2 => \N__44450\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40082\,
            in2 => \N__40013\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39890\,
            in2 => \N__39956\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44219\,
            in2 => \N__44153\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38402\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44623\,
            in2 => \N__44648\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40457\,
            in2 => \N__40488\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40379\,
            in2 => \N__46590\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46430\,
            in2 => \N__38525\,
            in3 => \N__38501\,
            lcout => \current_shift_inst.un38_control_input_0_s1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40526\,
            in2 => \N__46591\,
            in3 => \N__38483\,
            lcout => \current_shift_inst.un38_control_input_0_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46434\,
            in2 => \N__40373\,
            in3 => \N__38465\,
            lcout => \current_shift_inst.un38_control_input_0_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40520\,
            in2 => \N__46592\,
            in3 => \N__38450\,
            lcout => \current_shift_inst.un38_control_input_0_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46438\,
            in2 => \N__40352\,
            in3 => \N__38432\,
            lcout => \current_shift_inst.un38_control_input_0_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46264\,
            in2 => \N__38924\,
            in3 => \N__38612\,
            lcout => \current_shift_inst.un38_control_input_0_s1_8\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40547\,
            in2 => \N__46442\,
            in3 => \N__38597\,
            lcout => \current_shift_inst.un38_control_input_0_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46268\,
            in2 => \N__41351\,
            in3 => \N__38582\,
            lcout => \current_shift_inst.un38_control_input_0_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40511\,
            in2 => \N__46443\,
            in3 => \N__38567\,
            lcout => \current_shift_inst.un38_control_input_0_s1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46272\,
            in2 => \N__41300\,
            in3 => \N__38552\,
            lcout => \current_shift_inst.un38_control_input_0_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40358\,
            in2 => \N__46444\,
            in3 => \N__38537\,
            lcout => \current_shift_inst.un38_control_input_0_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46276\,
            in2 => \N__41636\,
            in3 => \N__38534\,
            lcout => \current_shift_inst.un38_control_input_0_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40364\,
            in2 => \N__46445\,
            in3 => \N__38531\,
            lcout => \current_shift_inst.un38_control_input_0_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46336\,
            in2 => \N__39131\,
            in3 => \N__38528\,
            lcout => \current_shift_inst.un38_control_input_0_s1_16\,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39185\,
            in2 => \N__46504\,
            in3 => \N__38741\,
            lcout => \current_shift_inst.un38_control_input_0_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46340\,
            in2 => \N__39089\,
            in3 => \N__38738\,
            lcout => \current_shift_inst.un38_control_input_0_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45350\,
            in2 => \N__46505\,
            in3 => \N__38720\,
            lcout => \current_shift_inst.un38_control_input_0_s1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46344\,
            in2 => \N__39314\,
            in3 => \N__38702\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45266\,
            in2 => \N__46506\,
            in3 => \N__38687\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46348\,
            in2 => \N__38987\,
            in3 => \N__38672\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41624\,
            in2 => \N__46507\,
            in3 => \N__38654\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38975\,
            in2 => \N__46508\,
            in3 => \N__38639\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46355\,
            in2 => \N__39116\,
            in3 => \N__38831\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41363\,
            in2 => \N__46509\,
            in3 => \N__38828\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46359\,
            in2 => \N__39101\,
            in3 => \N__38825\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39323\,
            in2 => \N__46510\,
            in3 => \N__38807\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46363\,
            in2 => \N__38966\,
            in3 => \N__38789\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40430\,
            in2 => \N__46511\,
            in3 => \N__38774\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__45999\,
            in1 => \N__46367\,
            in2 => \_gnd_net_\,
            in3 => \N__38771\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45986\,
            in1 => \N__47140\,
            in2 => \N__46623\,
            in3 => \N__44598\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__46041\,
            in1 => \N__46524\,
            in2 => \N__47056\,
            in3 => \N__45987\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45984\,
            in1 => \N__46735\,
            in2 => \N__46622\,
            in3 => \N__40732\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47049\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \N__46525\,
            in1 => \N__45408\,
            in2 => \N__46009\,
            in3 => \N__47012\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__47256\,
            in1 => \N__45985\,
            in2 => \N__46700\,
            in3 => \N__46523\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47255\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46781\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__41823\,
            in1 => \N__38912\,
            in2 => \_gnd_net_\,
            in3 => \N__38903\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38885\,
            in1 => \N__38876\,
            in2 => \_gnd_net_\,
            in3 => \N__41822\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__41826\,
            in1 => \N__38858\,
            in2 => \_gnd_net_\,
            in3 => \N__38849\,
            lcout => \current_shift_inst.control_input_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__39074\,
            in1 => \N__39068\,
            in2 => \_gnd_net_\,
            in3 => \N__41824\,
            lcout => \current_shift_inst.control_input_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__41825\,
            in1 => \N__39050\,
            in2 => \_gnd_net_\,
            in3 => \N__39044\,
            lcout => \current_shift_inst.control_input_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__41827\,
            in1 => \N__39023\,
            in2 => \_gnd_net_\,
            in3 => \N__39014\,
            lcout => \current_shift_inst.control_input_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45994\,
            in1 => \N__46527\,
            in2 => \N__47516\,
            in3 => \N__45367\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46526\,
            in1 => \N__45995\,
            in2 => \N__47432\,
            in3 => \N__45285\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46625\,
            in1 => \N__45882\,
            in2 => \N__47384\,
            in3 => \N__42178\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45883\,
            in1 => \N__46627\,
            in2 => \N__48055\,
            in3 => \N__42052\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46626\,
            in1 => \N__45887\,
            in2 => \N__47836\,
            in3 => \N__41982\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45885\,
            in1 => \N__46630\,
            in2 => \N__47969\,
            in3 => \N__42021\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46628\,
            in1 => \N__45884\,
            in2 => \N__48014\,
            in3 => \N__42080\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45881\,
            in1 => \N__46629\,
            in2 => \N__47600\,
            in3 => \N__45630\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46624\,
            in1 => \N__45886\,
            in2 => \N__47924\,
            in3 => \N__41948\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__39167\,
            in1 => \N__39158\,
            in2 => \_gnd_net_\,
            in3 => \N__41862\,
            lcout => \current_shift_inst.control_input_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46637\,
            in1 => \N__46008\,
            in2 => \N__47840\,
            in3 => \N__41983\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__45249\,
            in1 => \N__46001\,
            in2 => \N__47648\,
            in3 => \N__46638\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46002\,
            in1 => \N__48010\,
            in2 => \N__46660\,
            in3 => \N__42079\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__46007\,
            in1 => \N__46632\,
            in2 => \N__47923\,
            in3 => \N__41947\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__46631\,
            in1 => \N__41917\,
            in2 => \N__47558\,
            in3 => \N__46005\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110011"
        )
    port map (
            in0 => \N__45029\,
            in1 => \N__46004\,
            in2 => \N__41012\,
            in3 => \N__46642\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46003\,
            in1 => \N__47875\,
            in2 => \N__46659\,
            in3 => \N__41716\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__46006\,
            in1 => \N__46636\,
            in2 => \N__47473\,
            in3 => \N__45465\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40000\,
            in1 => \N__44059\,
            in2 => \_gnd_net_\,
            in3 => \N__50398\,
            lcout => \elapsed_time_ns_1_RNI47DN9_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39292\,
            in1 => \N__42630\,
            in2 => \_gnd_net_\,
            in3 => \N__50397\,
            lcout => \elapsed_time_ns_1_RNIG23T9_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_16_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__39542\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39256\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_16_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__39541\,
            in1 => \N__39272\,
            in2 => \_gnd_net_\,
            in3 => \N__39255\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39232\,
            in1 => \N__42666\,
            in2 => \_gnd_net_\,
            in3 => \N__50399\,
            lcout => \elapsed_time_ns_1_RNIF13T9_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39438\,
            in2 => \_gnd_net_\,
            in3 => \N__39469\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39571\,
            in1 => \N__43702\,
            in2 => \_gnd_net_\,
            in3 => \N__50400\,
            lcout => \elapsed_time_ns_1_RNIE03T9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39550\,
            in2 => \_gnd_net_\,
            in3 => \N__39506\,
            lcout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39458\,
            in3 => \N__39437\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__39398\,
            in1 => \N__39376\,
            in2 => \N__39344\,
            in3 => \N__39689\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50405\,
            in1 => \N__40215\,
            in2 => \_gnd_net_\,
            in3 => \N__42450\,
            lcout => \elapsed_time_ns_1_RNIJ53T9_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__39688\,
            in1 => \N__39397\,
            in2 => \N__39380\,
            in3 => \N__39340\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43840\,
            in1 => \N__39874\,
            in2 => \_gnd_net_\,
            in3 => \N__50407\,
            lcout => \elapsed_time_ns_1_RNI7ADN9_0_29\,
            ltout => \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_29_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50409\,
            in1 => \_gnd_net_\,
            in2 => \N__39347\,
            in3 => \N__43841\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50037\,
            ce => \N__49566\,
            sr => \N__49096\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43912\,
            in1 => \N__39967\,
            in2 => \_gnd_net_\,
            in3 => \N__50406\,
            lcout => \elapsed_time_ns_1_RNI69DN9_0_28\,
            ltout => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_28_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50408\,
            in1 => \_gnd_net_\,
            in2 => \N__39692\,
            in3 => \N__43913\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50037\,
            ce => \N__49566\,
            sr => \N__49096\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__39667\,
            in1 => \N__39648\,
            in2 => \N__39614\,
            in3 => \N__39599\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__39598\,
            in1 => \N__39666\,
            in2 => \N__39653\,
            in3 => \N__39610\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43251\,
            in1 => \N__40417\,
            in2 => \_gnd_net_\,
            in3 => \N__50291\,
            lcout => \elapsed_time_ns_1_RNI14DN9_0_23\,
            ltout => \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_23_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50293\,
            in1 => \_gnd_net_\,
            in2 => \N__39617\,
            in3 => \N__43252\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50030\,
            ce => \N__49460\,
            sr => \N__49102\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43308\,
            in1 => \N__40114\,
            in2 => \_gnd_net_\,
            in3 => \N__50290\,
            lcout => \elapsed_time_ns_1_RNI03DN9_0_22\,
            ltout => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_22_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50292\,
            in1 => \_gnd_net_\,
            in2 => \N__39602\,
            in3 => \N__43309\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50030\,
            ce => \N__49460\,
            sr => \N__49102\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__39845\,
            in1 => \N__39835\,
            in2 => \N__50074\,
            in3 => \N__39820\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50556\,
            in1 => \N__50590\,
            in2 => \_gnd_net_\,
            in3 => \N__50281\,
            lcout => \elapsed_time_ns_1_RNI04EN9_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__41183\,
            in1 => \N__41024\,
            in2 => \N__41141\,
            in3 => \N__50589\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44140\,
            in2 => \N__39851\,
            in3 => \N__44101\,
            lcout => \elapsed_time_ns_1_RNIV2EN9_0_30\,
            ltout => \elapsed_time_ns_1_RNIV2EN9_0_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_30_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__44141\,
            in1 => \_gnd_net_\,
            in2 => \N__39848\,
            in3 => \N__50283\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50017\,
            ce => \N__49520\,
            sr => \N__49107\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__39844\,
            in1 => \N__39834\,
            in2 => \N__50075\,
            in3 => \N__39819\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41120\,
            in1 => \N__42977\,
            in2 => \_gnd_net_\,
            in3 => \N__50282\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50017\,
            ce => \N__49520\,
            sr => \N__49107\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__39772\,
            in1 => \N__39751\,
            in2 => \N__39704\,
            in3 => \N__39713\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__39712\,
            in1 => \N__39773\,
            in2 => \N__39752\,
            in3 => \N__39700\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40868\,
            in1 => \N__42812\,
            in2 => \_gnd_net_\,
            in3 => \N__50327\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50007\,
            ce => \N__45118\,
            sr => \N__49112\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50325\,
            in1 => \N__42743\,
            in2 => \_gnd_net_\,
            in3 => \N__40901\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50007\,
            ce => \N__45118\,
            sr => \N__49112\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40843\,
            in1 => \N__42932\,
            in2 => \_gnd_net_\,
            in3 => \N__50326\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50007\,
            ce => \N__45118\,
            sr => \N__49112\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__40070\,
            in1 => \N__40045\,
            in2 => \N__40037\,
            in3 => \N__39980\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__39979\,
            in1 => \N__40069\,
            in2 => \N__40049\,
            in3 => \N__40036\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_26_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40001\,
            in1 => \N__44058\,
            in2 => \_gnd_net_\,
            in3 => \N__50511\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49997\,
            ce => \N__45116\,
            sr => \N__49119\
        );

    \phase_controller_inst2.stoper_hc.target_time_28_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43911\,
            in1 => \N__39971\,
            in2 => \_gnd_net_\,
            in3 => \N__50512\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49997\,
            ce => \N__45116\,
            sr => \N__49119\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__39898\,
            in1 => \N__39944\,
            in2 => \N__39923\,
            in3 => \N__39859\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__39943\,
            in1 => \N__39919\,
            in2 => \N__39863\,
            in3 => \N__39899\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_29_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50510\,
            in1 => \N__43839\,
            in2 => \_gnd_net_\,
            in3 => \N__39878\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49997\,
            ce => \N__45116\,
            sr => \N__49119\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__40334\,
            in1 => \N__40309\,
            in2 => \N__40229\,
            in3 => \N__40265\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__40264\,
            in1 => \N__40333\,
            in2 => \N__40313\,
            in3 => \N__40225\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_20_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43427\,
            in1 => \N__40283\,
            in2 => \_gnd_net_\,
            in3 => \N__50354\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49986\,
            ce => \N__45113\,
            sr => \N__49126\
        );

    \phase_controller_inst2.stoper_hc.target_time_21_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50351\,
            in1 => \N__40256\,
            in2 => \_gnd_net_\,
            in3 => \N__43370\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49986\,
            ce => \N__45113\,
            sr => \N__49126\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__40217\,
            in1 => \N__50353\,
            in2 => \_gnd_net_\,
            in3 => \N__42454\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49986\,
            ce => \N__45113\,
            sr => \N__49126\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50352\,
            in1 => \N__41063\,
            in2 => \_gnd_net_\,
            in3 => \N__42326\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49986\,
            ce => \N__45113\,
            sr => \N__49126\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__40406\,
            in1 => \N__40103\,
            in2 => \N__40169\,
            in3 => \N__40146\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__40102\,
            in1 => \N__40168\,
            in2 => \N__40148\,
            in3 => \N__40405\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_22_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43313\,
            in1 => \N__40121\,
            in2 => \_gnd_net_\,
            in3 => \N__50509\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49976\,
            ce => \N__45111\,
            sr => \N__49132\
        );

    \phase_controller_inst2.stoper_hc.target_time_23_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50507\,
            in1 => \N__43253\,
            in2 => \_gnd_net_\,
            in3 => \N__40421\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49976\,
            ce => \N__45111\,
            sr => \N__49132\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50505\,
            in1 => \N__41174\,
            in2 => \_gnd_net_\,
            in3 => \N__43085\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49976\,
            ce => \N__45111\,
            sr => \N__49132\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43157\,
            in1 => \N__41096\,
            in2 => \_gnd_net_\,
            in3 => \N__50508\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49976\,
            ce => \N__45111\,
            sr => \N__49132\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50506\,
            in1 => \N__42710\,
            in2 => \_gnd_net_\,
            in3 => \N__43028\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49976\,
            ce => \N__45111\,
            sr => \N__49132\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45911\,
            in1 => \N__46650\,
            in2 => \N__46931\,
            in3 => \N__40609\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46644\,
            in1 => \N__45913\,
            in2 => \N__46793\,
            in3 => \N__44551\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45918\,
            in1 => \N__46649\,
            in2 => \N__45215\,
            in3 => \N__47689\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46648\,
            in1 => \N__45917\,
            in2 => \N__47060\,
            in3 => \N__46045\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45915\,
            in1 => \N__46646\,
            in2 => \N__40709\,
            in3 => \N__47306\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46643\,
            in1 => \N__45912\,
            in2 => \N__46840\,
            in3 => \N__41338\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45914\,
            in1 => \N__46645\,
            in2 => \N__40736\,
            in3 => \N__46736\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46647\,
            in1 => \N__45916\,
            in2 => \N__47144\,
            in3 => \N__44605\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__40489\,
            in1 => \N__40627\,
            in2 => \N__40451\,
            in3 => \N__45826\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48296\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49963\,
            ce => \N__47794\,
            sr => \N__49145\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40445\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110100011"
        )
    port map (
            in0 => \N__40628\,
            in1 => \N__40450\,
            in2 => \N__45910\,
            in3 => \N__40490\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__45519\,
            in1 => \N__40626\,
            in2 => \_gnd_net_\,
            in3 => \N__40446\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \N__46601\,
            in1 => \N__45830\,
            in2 => \N__45028\,
            in3 => \N__41008\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__47218\,
            in1 => \N__45991\,
            in2 => \N__40667\,
            in3 => \N__46513\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45992\,
            in1 => \N__47219\,
            in2 => \N__46621\,
            in3 => \N__40666\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45993\,
            in2 => \_gnd_net_\,
            in3 => \N__46512\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47217\,
            in1 => \N__45518\,
            in2 => \_gnd_net_\,
            in3 => \N__40662\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45671\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__45672\,
            in1 => \_gnd_net_\,
            in2 => \N__40529\,
            in3 => \N__45517\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47762\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49954\,
            ce => \N__47793\,
            sr => \N__49152\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47726\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49954\,
            ce => \N__47793\,
            sr => \N__49152\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45521\,
            in1 => \N__46867\,
            in2 => \_gnd_net_\,
            in3 => \N__40573\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46827\,
            in1 => \N__45522\,
            in2 => \_gnd_net_\,
            in3 => \N__41331\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45525\,
            in1 => \N__47301\,
            in2 => \_gnd_net_\,
            in3 => \N__40695\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46917\,
            in1 => \N__45520\,
            in2 => \_gnd_net_\,
            in3 => \N__40602\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45526\,
            in1 => \N__47260\,
            in2 => \_gnd_net_\,
            in3 => \N__46686\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46731\,
            in1 => \N__45524\,
            in2 => \_gnd_net_\,
            in3 => \N__40728\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45523\,
            in1 => \N__46782\,
            in2 => \_gnd_net_\,
            in3 => \N__44541\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47431\,
            in1 => \N__45527\,
            in2 => \_gnd_net_\,
            in3 => \N__45286\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40637\,
            in2 => \N__45085\,
            in3 => \N__45081\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41957\,
            in2 => \_gnd_net_\,
            in3 => \N__40586\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42149\,
            in3 => \N__40562\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45602\,
            in2 => \_gnd_net_\,
            in3 => \N__40748\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40745\,
            in2 => \_gnd_net_\,
            in3 => \N__40739\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46970\,
            in2 => \_gnd_net_\,
            in3 => \N__40712\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45437\,
            in2 => \_gnd_net_\,
            in3 => \N__40679\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40676\,
            in2 => \_gnd_net_\,
            in3 => \N__40670\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46940\,
            in2 => \_gnd_net_\,
            in3 => \N__40649\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_16_18_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41990\,
            in2 => \_gnd_net_\,
            in3 => \N__40646\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44564\,
            in2 => \_gnd_net_\,
            in3 => \N__40643\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42107\,
            in2 => \_gnd_net_\,
            in3 => \N__40640\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40781\,
            in2 => \_gnd_net_\,
            in3 => \N__40775\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46949\,
            in2 => \_gnd_net_\,
            in3 => \N__40772\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46958\,
            in2 => \_gnd_net_\,
            in3 => \N__40769\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42260\,
            in2 => \_gnd_net_\,
            in3 => \N__40766\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42137\,
            in2 => \_gnd_net_\,
            in3 => \N__40763\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42245\,
            in2 => \_gnd_net_\,
            in3 => \N__40760\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42227\,
            in2 => \_gnd_net_\,
            in3 => \N__40757\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42131\,
            in3 => \N__40754\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42098\,
            in2 => \_gnd_net_\,
            in3 => \N__40751\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42113\,
            in2 => \_gnd_net_\,
            in3 => \N__40808\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42089\,
            in2 => \_gnd_net_\,
            in3 => \N__40805\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42236\,
            in2 => \_gnd_net_\,
            in3 => \N__40802\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42266\,
            in2 => \_gnd_net_\,
            in3 => \N__40799\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_16_20_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42206\,
            in2 => \_gnd_net_\,
            in3 => \N__40796\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42251\,
            in2 => \_gnd_net_\,
            in3 => \N__40793\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42215\,
            in2 => \_gnd_net_\,
            in3 => \N__40790\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42197\,
            in3 => \N__40787\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40784\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46000\,
            in2 => \_gnd_net_\,
            in3 => \N__41001\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_17_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40860\,
            in1 => \N__42811\,
            in2 => \_gnd_net_\,
            in3 => \N__50501\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50050\,
            ce => \N__49550\,
            sr => \N__49088\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__40973\,
            in1 => \N__40961\,
            in2 => \N__40880\,
            in3 => \N__40936\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__40972\,
            in1 => \N__40960\,
            in2 => \N__40937\,
            in3 => \N__40876\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42741\,
            in1 => \N__40894\,
            in2 => \_gnd_net_\,
            in3 => \N__50403\,
            lcout => \elapsed_time_ns_1_RNI46CN9_0_17\,
            ltout => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50404\,
            in1 => \_gnd_net_\,
            in2 => \N__40883\,
            in3 => \N__42742\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50047\,
            ce => \N__49544\,
            sr => \N__49089\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42804\,
            in1 => \N__40864\,
            in2 => \_gnd_net_\,
            in3 => \N__50402\,
            lcout => \elapsed_time_ns_1_RNI35CN9_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_17_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50401\,
            in1 => \N__40836\,
            in2 => \_gnd_net_\,
            in3 => \N__42927\,
            lcout => \elapsed_time_ns_1_RNI13CN9_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40844\,
            in1 => \N__42928\,
            in2 => \_gnd_net_\,
            in3 => \N__50410\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50043\,
            ce => \N__49501\,
            sr => \N__49093\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41055\,
            in1 => \N__42322\,
            in2 => \_gnd_net_\,
            in3 => \N__50411\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50043\,
            ce => \N__49501\,
            sr => \N__49093\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43145\,
            in1 => \N__41089\,
            in2 => \_gnd_net_\,
            in3 => \N__50294\,
            lcout => \elapsed_time_ns_1_RNITUBN9_0_10\,
            ltout => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50296\,
            in1 => \_gnd_net_\,
            in2 => \N__41078\,
            in3 => \N__43146\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50038\,
            ce => \N__49563\,
            sr => \N__49097\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50295\,
            in1 => \N__41059\,
            in2 => \_gnd_net_\,
            in3 => \N__42318\,
            lcout => \elapsed_time_ns_1_RNIL73T9_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50297\,
            in1 => \N__41166\,
            in2 => \_gnd_net_\,
            in3 => \N__43078\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50038\,
            ce => \N__49563\,
            sr => \N__49097\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42363\,
            in2 => \_gnd_net_\,
            in3 => \N__42432\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44505\,
            in1 => \N__42612\,
            in2 => \N__43700\,
            in3 => \N__42648\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43968\,
            in2 => \N__41027\,
            in3 => \N__43905\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43076\,
            in1 => \N__42317\,
            in2 => \N__43150\,
            in3 => \N__43016\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__42556\,
            in1 => \N__42503\,
            in2 => \N__41192\,
            in3 => \N__41189\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43077\,
            in1 => \N__41170\,
            in2 => \_gnd_net_\,
            in3 => \N__50298\,
            lcout => \elapsed_time_ns_1_RNIUVBN9_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__43017\,
            in1 => \_gnd_net_\,
            in2 => \N__50420\,
            in3 => \N__42709\,
            lcout => \elapsed_time_ns_1_RNIV0CN9_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43476\,
            in1 => \N__43544\,
            in2 => \N__43416\,
            in3 => \N__42726\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42858\,
            in1 => \N__42917\,
            in2 => \N__42803\,
            in3 => \N__42971\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41126\,
            in1 => \N__41132\,
            in2 => \N__41150\,
            in3 => \N__41147\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44364\,
            in1 => \N__43236\,
            in2 => \N__43299\,
            in3 => \N__43350\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44139\,
            in1 => \N__44037\,
            in2 => \N__44256\,
            in3 => \N__43827\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42972\,
            in1 => \N__41119\,
            in2 => \_gnd_net_\,
            in3 => \N__50302\,
            lcout => \elapsed_time_ns_1_RNI02CN9_0_13\,
            ltout => \elapsed_time_ns_1_RNI02CN9_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50303\,
            in1 => \_gnd_net_\,
            in2 => \N__41231\,
            in3 => \N__42973\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50018\,
            ce => \N__45119\,
            sr => \N__49108\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41535\,
            in1 => \N__43749\,
            in2 => \_gnd_net_\,
            in3 => \N__41216\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__50008\,
            ce => \N__41432\,
            sr => \N__49113\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41541\,
            in1 => \N__43722\,
            in2 => \_gnd_net_\,
            in3 => \N__41213\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__50008\,
            ce => \N__41432\,
            sr => \N__49113\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41536\,
            in1 => \N__42594\,
            in2 => \_gnd_net_\,
            in3 => \N__41210\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__50008\,
            ce => \N__41432\,
            sr => \N__49113\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41542\,
            in1 => \N__42540\,
            in2 => \_gnd_net_\,
            in3 => \N__41207\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__50008\,
            ce => \N__41432\,
            sr => \N__49113\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41537\,
            in1 => \N__42471\,
            in2 => \_gnd_net_\,
            in3 => \N__41204\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__50008\,
            ce => \N__41432\,
            sr => \N__49113\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41543\,
            in1 => \N__42405\,
            in2 => \_gnd_net_\,
            in3 => \N__41201\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__50008\,
            ce => \N__41432\,
            sr => \N__49113\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41538\,
            in1 => \N__42340\,
            in2 => \_gnd_net_\,
            in3 => \N__41198\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__50008\,
            ce => \N__41432\,
            sr => \N__49113\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41544\,
            in1 => \N__42282\,
            in2 => \_gnd_net_\,
            in3 => \N__41195\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__50008\,
            ce => \N__41432\,
            sr => \N__49113\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41560\,
            in1 => \N__43107\,
            in2 => \_gnd_net_\,
            in3 => \N__41258\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__49998\,
            ce => \N__41431\,
            sr => \N__49120\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41548\,
            in1 => \N__43047\,
            in2 => \_gnd_net_\,
            in3 => \N__41255\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__49998\,
            ce => \N__41431\,
            sr => \N__49120\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41557\,
            in1 => \N__42993\,
            in2 => \_gnd_net_\,
            in3 => \N__41252\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__49998\,
            ce => \N__41431\,
            sr => \N__49120\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41545\,
            in1 => \N__42948\,
            in2 => \_gnd_net_\,
            in3 => \N__41249\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__49998\,
            ce => \N__41431\,
            sr => \N__49120\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41558\,
            in1 => \N__42888\,
            in2 => \_gnd_net_\,
            in3 => \N__41246\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__49998\,
            ce => \N__41431\,
            sr => \N__49120\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41546\,
            in1 => \N__42826\,
            in2 => \_gnd_net_\,
            in3 => \N__41243\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__49998\,
            ce => \N__41431\,
            sr => \N__49120\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41559\,
            in1 => \N__42759\,
            in2 => \_gnd_net_\,
            in3 => \N__41240\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__49998\,
            ce => \N__41431\,
            sr => \N__49120\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41547\,
            in1 => \N__43573\,
            in2 => \_gnd_net_\,
            in3 => \N__41237\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__49998\,
            ce => \N__41431\,
            sr => \N__49120\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41549\,
            in1 => \N__43512\,
            in2 => \_gnd_net_\,
            in3 => \N__41234\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__49987\,
            ce => \N__41430\,
            sr => \N__49127\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41561\,
            in1 => \N__43449\,
            in2 => \_gnd_net_\,
            in3 => \N__41285\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__49987\,
            ce => \N__41430\,
            sr => \N__49127\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41550\,
            in1 => \N__43386\,
            in2 => \_gnd_net_\,
            in3 => \N__41282\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__49987\,
            ce => \N__41430\,
            sr => \N__49127\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41562\,
            in1 => \N__43329\,
            in2 => \_gnd_net_\,
            in3 => \N__41279\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__49987\,
            ce => \N__41430\,
            sr => \N__49127\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41551\,
            in1 => \N__43269\,
            in2 => \_gnd_net_\,
            in3 => \N__41276\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__49987\,
            ce => \N__41430\,
            sr => \N__49127\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41563\,
            in1 => \N__43204\,
            in2 => \_gnd_net_\,
            in3 => \N__41273\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__49987\,
            ce => \N__41430\,
            sr => \N__49127\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41552\,
            in1 => \N__43176\,
            in2 => \_gnd_net_\,
            in3 => \N__41270\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__49987\,
            ce => \N__41430\,
            sr => \N__49127\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41564\,
            in1 => \N__44079\,
            in2 => \_gnd_net_\,
            in3 => \N__41267\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__49987\,
            ce => \N__41430\,
            sr => \N__49127\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41553\,
            in1 => \N__44007\,
            in2 => \_gnd_net_\,
            in3 => \N__41264\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__49977\,
            ce => \N__41420\,
            sr => \N__49133\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41539\,
            in1 => \N__43935\,
            in2 => \_gnd_net_\,
            in3 => \N__41261\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__49977\,
            ce => \N__41420\,
            sr => \N__49133\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41554\,
            in1 => \N__43875\,
            in2 => \_gnd_net_\,
            in3 => \N__41573\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__49977\,
            ce => \N__41420\,
            sr => \N__49133\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41540\,
            in1 => \N__43779\,
            in2 => \_gnd_net_\,
            in3 => \N__41570\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__49977\,
            ce => \N__41420\,
            sr => \N__49133\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41555\,
            in1 => \N__43855\,
            in2 => \_gnd_net_\,
            in3 => \N__41567\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__49977\,
            ce => \N__41420\,
            sr => \N__49133\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__43804\,
            in1 => \N__41556\,
            in2 => \_gnd_net_\,
            in3 => \N__41435\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49977\,
            ce => \N__41420\,
            sr => \N__49133\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45838\,
            in1 => \N__46610\,
            in2 => \N__45257\,
            in3 => \N__47644\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45909\,
            in1 => \N__47968\,
            in2 => \N__46653\,
            in3 => \N__42026\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45835\,
            in1 => \N__46603\,
            in2 => \N__47186\,
            in3 => \N__46094\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46602\,
            in1 => \N__45834\,
            in2 => \N__46841\,
            in3 => \N__41339\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__47098\,
            in1 => \N__45907\,
            in2 => \N__45332\,
            in3 => \N__46605\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46604\,
            in1 => \N__45836\,
            in2 => \N__47102\,
            in3 => \N__45331\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__45837\,
            in1 => \N__47011\,
            in2 => \N__45419\,
            in3 => \N__46606\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45908\,
            in1 => \N__47341\,
            in2 => \N__46652\,
            in3 => \N__45169\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45003\,
            in2 => \N__45055\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44973\,
            in2 => \N__41612\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41603\,
            in2 => \N__44988\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44977\,
            in2 => \N__41597\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41588\,
            in2 => \N__44989\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44981\,
            in2 => \N__41582\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41684\,
            in2 => \N__44990\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44985\,
            in2 => \N__41678\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44937\,
            in2 => \N__41669\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44961\,
            in2 => \N__41660\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44934\,
            in2 => \N__45341\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44958\,
            in2 => \N__44579\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44935\,
            in2 => \N__45302\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44959\,
            in2 => \N__46019\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44936\,
            in2 => \N__45383\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44960\,
            in2 => \N__45428\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44918\,
            in2 => \N__45224\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45608\,
            in2 => \N__44969\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44922\,
            in2 => \N__41900\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42122\,
            in2 => \N__44970\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44926\,
            in2 => \N__45446\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41690\,
            in2 => \N__44971\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44930\,
            in2 => \N__42161\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45134\,
            in2 => \N__44972\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44905\,
            in2 => \N__42035\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42062\,
            in2 => \N__44966\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44909\,
            in2 => \N__41999\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41930\,
            in2 => \N__44967\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44913\,
            in2 => \N__41699\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41963\,
            in2 => \N__44968\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44917\,
            in2 => \N__41888\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__46010\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41876\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47868\,
            in1 => \N__45870\,
            in2 => \_gnd_net_\,
            in3 => \N__41715\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45869\,
            in1 => \N__48003\,
            in2 => \_gnd_net_\,
            in3 => \N__42078\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48042\,
            in1 => \N__45588\,
            in2 => \_gnd_net_\,
            in3 => \N__42051\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__47955\,
            in1 => \N__45872\,
            in2 => \N__42022\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47163\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45871\,
            in1 => \_gnd_net_\,
            in2 => \N__41984\,
            in3 => \N__47823\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46904\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47910\,
            in1 => \N__45873\,
            in2 => \_gnd_net_\,
            in3 => \N__41946\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45585\,
            in1 => \N__47541\,
            in2 => \_gnd_net_\,
            in3 => \N__41916\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47367\,
            in1 => \N__45586\,
            in2 => \_gnd_net_\,
            in3 => \N__42177\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46855\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47577\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47446\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45587\,
            in1 => \N__47494\,
            in2 => \_gnd_net_\,
            in3 => \N__45366\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47366\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47090\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47408\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47322\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47993\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47624\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47900\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47540\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48033\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47493\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47859\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47945\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47814\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_18_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42705\,
            in1 => \N__43024\,
            in2 => \_gnd_net_\,
            in3 => \N__50521\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50048\,
            ce => \N__49564\,
            sr => \N__49090\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42595\,
            in2 => \N__43757\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_18_7_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__50044\,
            ce => \N__43652\,
            sr => \N__49094\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42541\,
            in2 => \N__43730\,
            in3 => \N__42599\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__50044\,
            ce => \N__43652\,
            sr => \N__49094\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42596\,
            in2 => \N__42478\,
            in3 => \N__42545\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__50044\,
            ce => \N__43652\,
            sr => \N__49094\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42542\,
            in2 => \N__42412\,
            in3 => \N__42482\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__50044\,
            ce => \N__43652\,
            sr => \N__49094\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42346\,
            in2 => \N__42479\,
            in3 => \N__42416\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__50044\,
            ce => \N__43652\,
            sr => \N__49094\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42289\,
            in2 => \N__42413\,
            in3 => \N__42350\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__50044\,
            ce => \N__43652\,
            sr => \N__49094\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42347\,
            in2 => \N__43120\,
            in3 => \N__42296\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__50044\,
            ce => \N__43652\,
            sr => \N__49094\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43054\,
            in2 => \N__42293\,
            in3 => \N__43124\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__50044\,
            ce => \N__43652\,
            sr => \N__49094\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42994\,
            in2 => \N__43121\,
            in3 => \N__43058\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_18_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__50039\,
            ce => \N__43651\,
            sr => \N__49098\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42949\,
            in2 => \N__43055\,
            in3 => \N__42998\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__50039\,
            ce => \N__43651\,
            sr => \N__49098\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42995\,
            in2 => \N__42895\,
            in3 => \N__42953\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__50039\,
            ce => \N__43651\,
            sr => \N__49098\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42950\,
            in2 => \N__42838\,
            in3 => \N__42899\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__50039\,
            ce => \N__43651\,
            sr => \N__49098\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42766\,
            in2 => \N__42896\,
            in3 => \N__42842\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__50039\,
            ce => \N__43651\,
            sr => \N__49098\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43579\,
            in2 => \N__42839\,
            in3 => \N__42773\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__50039\,
            ce => \N__43651\,
            sr => \N__49098\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43519\,
            in2 => \N__42770\,
            in3 => \N__42713\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__50039\,
            ce => \N__43651\,
            sr => \N__49098\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43580\,
            in2 => \N__43460\,
            in3 => \N__43526\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__50039\,
            ce => \N__43651\,
            sr => \N__49098\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43387\,
            in2 => \N__43523\,
            in3 => \N__43463\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_18_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__50031\,
            ce => \N__43650\,
            sr => \N__49103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43330\,
            in2 => \N__43459\,
            in3 => \N__43391\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__50031\,
            ce => \N__43650\,
            sr => \N__49103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43388\,
            in2 => \N__43276\,
            in3 => \N__43334\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__50031\,
            ce => \N__43650\,
            sr => \N__49103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43331\,
            in2 => \N__43216\,
            in3 => \N__43280\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__50031\,
            ce => \N__43650\,
            sr => \N__49103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43183\,
            in2 => \N__43277\,
            in3 => \N__43220\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__50031\,
            ce => \N__43650\,
            sr => \N__49103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44086\,
            in2 => \N__43217\,
            in3 => \N__43190\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__50031\,
            ce => \N__43650\,
            sr => \N__49103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44014\,
            in2 => \N__43187\,
            in3 => \N__43160\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__50031\,
            ce => \N__43650\,
            sr => \N__49103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43942\,
            in2 => \N__44090\,
            in3 => \N__44021\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__50031\,
            ce => \N__43650\,
            sr => \N__49103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43876\,
            in2 => \N__44018\,
            in3 => \N__43946\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_18_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__50019\,
            ce => \N__43649\,
            sr => \N__49109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43786\,
            in2 => \N__43943\,
            in3 => \N__43880\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__50019\,
            ce => \N__43649\,
            sr => \N__49109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43877\,
            in2 => \N__43859\,
            in3 => \N__43811\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__50019\,
            ce => \N__43649\,
            sr => \N__49109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43808\,
            in2 => \N__43790\,
            in3 => \N__43763\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__50019\,
            ce => \N__43649\,
            sr => \N__49109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43760\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50019\,
            ce => \N__43649\,
            sr => \N__49109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43750\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50009\,
            ce => \N__43645\,
            sr => \N__49114\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43723\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50009\,
            ce => \N__43645\,
            sr => \N__49114\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44466\,
            in1 => \N__44499\,
            in2 => \_gnd_net_\,
            in3 => \N__50469\,
            lcout => \elapsed_time_ns_1_RNIDV2T9_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__44437\,
            in1 => \N__44416\,
            in2 => \N__44231\,
            in3 => \N__44321\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__44320\,
            in1 => \N__44438\,
            in2 => \N__44420\,
            in3 => \N__44227\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_24_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44385\,
            in1 => \N__44351\,
            in2 => \_gnd_net_\,
            in3 => \N__50514\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49999\,
            ce => \N__45117\,
            sr => \N__49121\
        );

    \phase_controller_inst2.stoper_hc.target_time_25_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50513\,
            in1 => \N__44312\,
            in2 => \_gnd_net_\,
            in3 => \N__44271\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49999\,
            ce => \N__45117\,
            sr => \N__49121\
        );

    \phase_controller_inst2.stoper_hc.target_time_31_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50588\,
            in1 => \N__50558\,
            in2 => \_gnd_net_\,
            in3 => \N__50515\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49999\,
            ce => \N__45117\,
            sr => \N__49121\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__45127\,
            in1 => \N__44200\,
            in2 => \N__44177\,
            in3 => \N__44209\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__44210\,
            in1 => \N__45128\,
            in2 => \N__44201\,
            in3 => \N__44176\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_30_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44138\,
            in1 => \N__44111\,
            in2 => \_gnd_net_\,
            in3 => \N__50528\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49988\,
            ce => \N__45114\,
            sr => \N__49128\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45086\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45813\,
            in2 => \N__45059\,
            in3 => \N__45685\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47757\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49978\,
            ce => \N__47795\,
            sr => \N__49134\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__45056\,
            in1 => \N__44986\,
            in2 => \_gnd_net_\,
            in3 => \N__45035\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__44987\,
            in1 => \_gnd_net_\,
            in2 => \N__44651\,
            in3 => \N__44641\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47130\,
            in1 => \N__45572\,
            in2 => \_gnd_net_\,
            in3 => \N__44606\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47129\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46587\,
            in1 => \N__45960\,
            in2 => \N__46789\,
            in3 => \N__44552\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47685\,
            in1 => \N__45552\,
            in2 => \_gnd_net_\,
            in3 => \N__45210\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__45551\,
            in1 => \N__47007\,
            in2 => \N__45415\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46589\,
            in1 => \N__45961\,
            in2 => \N__47512\,
            in3 => \N__45374\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47179\,
            in1 => \N__45549\,
            in2 => \_gnd_net_\,
            in3 => \N__46092\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45550\,
            in1 => \N__47091\,
            in2 => \_gnd_net_\,
            in3 => \N__45327\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45962\,
            in1 => \N__46588\,
            in2 => \N__45293\,
            in3 => \N__47421\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47643\,
            in1 => \N__45590\,
            in2 => \_gnd_net_\,
            in3 => \N__45250\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45959\,
            in1 => \N__46658\,
            in2 => \N__47690\,
            in3 => \N__45211\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47340\,
            in1 => \N__45591\,
            in2 => \_gnd_net_\,
            in3 => \N__45168\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45957\,
            in1 => \N__46657\,
            in2 => \N__47261\,
            in3 => \N__46699\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47178\,
            in1 => \N__45958\,
            in2 => \N__46661\,
            in3 => \N__46093\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47048\,
            in1 => \N__45589\,
            in2 => \_gnd_net_\,
            in3 => \N__46046\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__45956\,
            in1 => \N__45695\,
            in2 => \_gnd_net_\,
            in3 => \N__45686\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45592\,
            in1 => \N__47595\,
            in2 => \_gnd_net_\,
            in3 => \N__45637\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46818\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45593\,
            in1 => \N__47460\,
            in2 => \_gnd_net_\,
            in3 => \N__45472\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47283\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46714\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47675\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47003\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47200\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48253\,
            in2 => \N__47722\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__49940\,
            ce => \N__47791\,
            sr => \N__49162\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48232\,
            in2 => \N__48292\,
            in3 => \N__46844\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__49940\,
            ce => \N__47791\,
            sr => \N__49162\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48254\,
            in2 => \N__48212\,
            in3 => \N__46796\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__49940\,
            ce => \N__47791\,
            sr => \N__49162\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48233\,
            in2 => \N__48182\,
            in3 => \N__46739\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__49940\,
            ce => \N__47791\,
            sr => \N__49162\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48211\,
            in2 => \N__48151\,
            in3 => \N__46703\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__49940\,
            ce => \N__47791\,
            sr => \N__49162\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48181\,
            in2 => \N__48121\,
            in3 => \N__47264\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__49940\,
            ce => \N__47791\,
            sr => \N__49162\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48088\,
            in2 => \N__48152\,
            in3 => \N__47222\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__49940\,
            ce => \N__47791\,
            sr => \N__49162\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48544\,
            in2 => \N__48122\,
            in3 => \N__47189\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__49940\,
            ce => \N__47791\,
            sr => \N__49162\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48517\,
            in2 => \N__48092\,
            in3 => \N__47147\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__49933\,
            ce => \N__47790\,
            sr => \N__49167\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48493\,
            in2 => \N__48548\,
            in3 => \N__47105\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__49933\,
            ce => \N__47790\,
            sr => \N__49167\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48518\,
            in2 => \N__48469\,
            in3 => \N__47063\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__49933\,
            ce => \N__47790\,
            sr => \N__49167\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48494\,
            in2 => \N__48439\,
            in3 => \N__47015\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__49933\,
            ce => \N__47790\,
            sr => \N__49167\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48409\,
            in2 => \N__48470\,
            in3 => \N__46973\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__49933\,
            ce => \N__47790\,
            sr => \N__49167\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48382\,
            in2 => \N__48440\,
            in3 => \N__47651\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__49933\,
            ce => \N__47790\,
            sr => \N__49167\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48410\,
            in2 => \N__48355\,
            in3 => \N__47603\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__49933\,
            ce => \N__47790\,
            sr => \N__49167\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48322\,
            in2 => \N__48386\,
            in3 => \N__47561\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__49933\,
            ce => \N__47790\,
            sr => \N__49167\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48760\,
            in2 => \N__48356\,
            in3 => \N__47519\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_18_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__49927\,
            ce => \N__47789\,
            sr => \N__49172\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48323\,
            in2 => \N__48739\,
            in3 => \N__47477\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__49927\,
            ce => \N__47789\,
            sr => \N__49172\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48761\,
            in2 => \N__48713\,
            in3 => \N__47435\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__49927\,
            ce => \N__47789\,
            sr => \N__49172\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48682\,
            in2 => \N__48740\,
            in3 => \N__47387\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__49927\,
            ce => \N__47789\,
            sr => \N__49172\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48712\,
            in2 => \N__48658\,
            in3 => \N__47348\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__49927\,
            ce => \N__47789\,
            sr => \N__49172\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48628\,
            in2 => \N__48686\,
            in3 => \N__48062\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__49927\,
            ce => \N__47789\,
            sr => \N__49172\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48604\,
            in2 => \N__48659\,
            in3 => \N__48017\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__49927\,
            ce => \N__47789\,
            sr => \N__49172\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48629\,
            in2 => \N__48578\,
            in3 => \N__47972\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__49927\,
            ce => \N__47789\,
            sr => \N__49172\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50851\,
            in2 => \N__48608\,
            in3 => \N__47927\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_18_22_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__49922\,
            ce => \N__47788\,
            sr => \N__49178\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48577\,
            in2 => \N__50827\,
            in3 => \N__47879\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__49922\,
            ce => \N__47788\,
            sr => \N__49178\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50801\,
            in2 => \N__50855\,
            in3 => \N__47843\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__49922\,
            ce => \N__47788\,
            sr => \N__49178\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50657\,
            in2 => \N__50828\,
            in3 => \N__47798\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__49922\,
            ce => \N__47788\,
            sr => \N__49178\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47765\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50758\,
            in1 => \N__47712\,
            in2 => \_gnd_net_\,
            in3 => \N__47693\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_23_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__49915\,
            ce => \N__50633\,
            sr => \N__49182\
        );

    \current_shift_inst.timer_s1.counter_1_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50754\,
            in1 => \N__48276\,
            in2 => \_gnd_net_\,
            in3 => \N__48257\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__49915\,
            ce => \N__50633\,
            sr => \N__49182\
        );

    \current_shift_inst.timer_s1.counter_2_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50759\,
            in1 => \N__48252\,
            in2 => \_gnd_net_\,
            in3 => \N__48236\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__49915\,
            ce => \N__50633\,
            sr => \N__49182\
        );

    \current_shift_inst.timer_s1.counter_3_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50755\,
            in1 => \N__48231\,
            in2 => \_gnd_net_\,
            in3 => \N__48215\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__49915\,
            ce => \N__50633\,
            sr => \N__49182\
        );

    \current_shift_inst.timer_s1.counter_4_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50760\,
            in1 => \N__48201\,
            in2 => \_gnd_net_\,
            in3 => \N__48185\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__49915\,
            ce => \N__50633\,
            sr => \N__49182\
        );

    \current_shift_inst.timer_s1.counter_5_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50756\,
            in1 => \N__48171\,
            in2 => \_gnd_net_\,
            in3 => \N__48155\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__49915\,
            ce => \N__50633\,
            sr => \N__49182\
        );

    \current_shift_inst.timer_s1.counter_6_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50761\,
            in1 => \N__48139\,
            in2 => \_gnd_net_\,
            in3 => \N__48125\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__49915\,
            ce => \N__50633\,
            sr => \N__49182\
        );

    \current_shift_inst.timer_s1.counter_7_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50757\,
            in1 => \N__48109\,
            in2 => \_gnd_net_\,
            in3 => \N__48095\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__49915\,
            ce => \N__50633\,
            sr => \N__49182\
        );

    \current_shift_inst.timer_s1.counter_8_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50779\,
            in1 => \N__48081\,
            in2 => \_gnd_net_\,
            in3 => \N__48065\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_24_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__49911\,
            ce => \N__50641\,
            sr => \N__49188\
        );

    \current_shift_inst.timer_s1.counter_9_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50783\,
            in1 => \N__48537\,
            in2 => \_gnd_net_\,
            in3 => \N__48521\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__49911\,
            ce => \N__50641\,
            sr => \N__49188\
        );

    \current_shift_inst.timer_s1.counter_10_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50776\,
            in1 => \N__48511\,
            in2 => \_gnd_net_\,
            in3 => \N__48497\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__49911\,
            ce => \N__50641\,
            sr => \N__49188\
        );

    \current_shift_inst.timer_s1.counter_11_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50780\,
            in1 => \N__48487\,
            in2 => \_gnd_net_\,
            in3 => \N__48473\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__49911\,
            ce => \N__50641\,
            sr => \N__49188\
        );

    \current_shift_inst.timer_s1.counter_12_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50777\,
            in1 => \N__48457\,
            in2 => \_gnd_net_\,
            in3 => \N__48443\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__49911\,
            ce => \N__50641\,
            sr => \N__49188\
        );

    \current_shift_inst.timer_s1.counter_13_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50781\,
            in1 => \N__48427\,
            in2 => \_gnd_net_\,
            in3 => \N__48413\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__49911\,
            ce => \N__50641\,
            sr => \N__49188\
        );

    \current_shift_inst.timer_s1.counter_14_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50778\,
            in1 => \N__48403\,
            in2 => \_gnd_net_\,
            in3 => \N__48389\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__49911\,
            ce => \N__50641\,
            sr => \N__49188\
        );

    \current_shift_inst.timer_s1.counter_15_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50782\,
            in1 => \N__48375\,
            in2 => \_gnd_net_\,
            in3 => \N__48359\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__49911\,
            ce => \N__50641\,
            sr => \N__49188\
        );

    \current_shift_inst.timer_s1.counter_16_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50762\,
            in1 => \N__48342\,
            in2 => \_gnd_net_\,
            in3 => \N__48326\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_18_25_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__49908\,
            ce => \N__50640\,
            sr => \N__49193\
        );

    \current_shift_inst.timer_s1.counter_17_LC_18_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50770\,
            in1 => \N__48315\,
            in2 => \_gnd_net_\,
            in3 => \N__48299\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__49908\,
            ce => \N__50640\,
            sr => \N__49193\
        );

    \current_shift_inst.timer_s1.counter_18_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50763\,
            in1 => \N__48759\,
            in2 => \_gnd_net_\,
            in3 => \N__48743\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__49908\,
            ce => \N__50640\,
            sr => \N__49193\
        );

    \current_shift_inst.timer_s1.counter_19_LC_18_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50771\,
            in1 => \N__48732\,
            in2 => \_gnd_net_\,
            in3 => \N__48716\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__49908\,
            ce => \N__50640\,
            sr => \N__49193\
        );

    \current_shift_inst.timer_s1.counter_20_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50764\,
            in1 => \N__48708\,
            in2 => \_gnd_net_\,
            in3 => \N__48689\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__49908\,
            ce => \N__50640\,
            sr => \N__49193\
        );

    \current_shift_inst.timer_s1.counter_21_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50772\,
            in1 => \N__48681\,
            in2 => \_gnd_net_\,
            in3 => \N__48662\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__49908\,
            ce => \N__50640\,
            sr => \N__49193\
        );

    \current_shift_inst.timer_s1.counter_22_LC_18_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50765\,
            in1 => \N__48646\,
            in2 => \_gnd_net_\,
            in3 => \N__48632\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__49908\,
            ce => \N__50640\,
            sr => \N__49193\
        );

    \current_shift_inst.timer_s1.counter_23_LC_18_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50773\,
            in1 => \N__48627\,
            in2 => \_gnd_net_\,
            in3 => \N__48611\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__49908\,
            ce => \N__50640\,
            sr => \N__49193\
        );

    \current_shift_inst.timer_s1.counter_24_LC_18_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50766\,
            in1 => \N__48597\,
            in2 => \_gnd_net_\,
            in3 => \N__48581\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_18_26_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__49905\,
            ce => \N__50642\,
            sr => \N__49199\
        );

    \current_shift_inst.timer_s1.counter_25_LC_18_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50774\,
            in1 => \N__48567\,
            in2 => \_gnd_net_\,
            in3 => \N__48551\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__49905\,
            ce => \N__50642\,
            sr => \N__49199\
        );

    \current_shift_inst.timer_s1.counter_26_LC_18_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50767\,
            in1 => \N__50850\,
            in2 => \_gnd_net_\,
            in3 => \N__50831\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__49905\,
            ce => \N__50642\,
            sr => \N__49199\
        );

    \current_shift_inst.timer_s1.counter_27_LC_18_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50775\,
            in1 => \N__50820\,
            in2 => \_gnd_net_\,
            in3 => \N__50804\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__49905\,
            ce => \N__50642\,
            sr => \N__49199\
        );

    \current_shift_inst.timer_s1.counter_28_LC_18_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50768\,
            in1 => \N__50800\,
            in2 => \_gnd_net_\,
            in3 => \N__50786\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__49905\,
            ce => \N__50642\,
            sr => \N__49199\
        );

    \current_shift_inst.timer_s1.counter_29_LC_18_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__50656\,
            in1 => \N__50769\,
            in2 => \_gnd_net_\,
            in3 => \N__50660\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49905\,
            ce => \N__50642\,
            sr => \N__49199\
        );

    \GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50054\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clock_output_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_31_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50591\,
            in1 => \N__50557\,
            in2 => \_gnd_net_\,
            in3 => \N__50524\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50045\,
            ce => \N__49542\,
            sr => \N__49104\
        );
end \INTERFACE\;
